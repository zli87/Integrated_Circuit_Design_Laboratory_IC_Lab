module INST_MEM_1 #(parameter ID_WIDTH=4, ADDR_WIDTH=32, DATA_WIDTH=16) (
// Glbal Signal
  	  input clk,
  	  input rst_n,
// slave interface
      // axi write address channel
      // src master
      input wire [ID_WIDTH-1:0]     awid_s_inf,
      input wire [ADDR_WIDTH-1:0] awaddr_s_inf,
      input wire [2:0]            awsize_s_inf,
      input wire [1:0]           awburst_s_inf,
      input wire [7:0]             awlen_s_inf,
      input wire                 awvalid_s_inf,
      // src slave
      output reg                 awready_s_inf,
      // -----------------------------

      // axi write data channel
      // src master
      input wire [DATA_WIDTH-1:0]  wdata_s_inf,
      input wire                   wlast_s_inf,
      input wire                  wvalid_s_inf,
      // src slave
      output reg                  wready_s_inf,

      // axi write response channel
      // src slave
      output reg  [ID_WIDTH-1:0]     bid_s_inf,
      output reg  [1:0]            bresp_s_inf,
      output reg                  bvalid_s_inf,
      // src master
      input wire                  bready_s_inf,
      // -----------------------------

      // axi read address channel
      // src master
      input wire [ID_WIDTH-1:0]     arid_s_inf,
      input wire [ADDR_WIDTH-1:0] araddr_s_inf,
      input wire [7:0]             arlen_s_inf,
      input wire [2:0]            arsize_s_inf,
      input wire [1:0]           arburst_s_inf,
      input wire                 arvalid_s_inf,
      // src slave
      output reg                 arready_s_inf,
      // -----------------------------

      // axi read data channel
      // slave
      output reg [ID_WIDTH-1:0]      rid_s_inf,
      output reg [DATA_WIDTH-1:0]  rdata_s_inf,
      output reg [1:0]             rresp_s_inf,
      output reg                   rlast_s_inf,
      output reg                  rvalid_s_inf,
      // master
      input wire                  rready_s_inf
      // -----------------------------
);
// Modify your "dat" in this directory path to initialized DRAM Value

parameter DRAM_p_r = "../00_TESTBED/DRAM/inst_1_file.dat";
// Modify DRAM_R_LAT           for Initial Read Data Latency,
//        DRAM_W_LAT           for Initial Write Data Latency
//        MAX_WAIT_READY_CYCLE for control the Upperlimit time to wait Response Ready Signal
//
//        reg [7:0] DRMA_r [0:8*1024-1] is the storage element in this simulation model

parameter DRAM_R_LAT = 90, DRAM_W_LAT =100, MAX_WAIT_READY_CYCLE=300;
reg	[7:0]	DRAM_r	[0:8*1024-1];

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Rstv0QmS+Pp9hT1xT+pSnfUdIDlFpjfaU9zziyHN5BaGTW6gIdFjx/TI9TxvpV0J
7SF6t1vU5bSAwOQrOylOizDnMl0dqoLnuPP17TMi3mgj9dSHpClAy2qDFdYosOm5
wjVXZMEmytoxurQWragZA4UueXCymOgkXb0mrE3QBTnU88RF0KXo9Q==
//pragma protect end_key_block
//pragma protect digest_block
oNzPyrjqSRmyc5ocNpjp494rV4k=
//pragma protect end_digest_block
//pragma protect data_block
idLlzWAVaA6wLPQxGLIdKSylzJinF+OO1MSNsQKwRzLmbZny0983PgsFfKJ8onz5
HcdTU5vLmc+Uf2wvykJdWtTJV8D53uwA4Pxw2pqo+llefrxRvzYA5S/93KmB0lne
xLCk61tmHQtlYVqwQDfd5e+VGYOv5Y1lsN8vXqwCepRsS6DB7+FEy4ikGrPNa7d6
UJ9/gRNb29K6r8Z+8q5g1EDbUXsGijWBqrwm84BZM1+0Vxr3pkun3yZCmo/CpG6n
2mX7vFmvh0cSSWWNBlk+EEP0g+zDVt9dP00A80Gsl+jzeu6JTuS0h6G2MhXDVLgg
1KbxAT07/dZkXtH2YgbP/5WjSP0fSqwqVRSN7l8nEqomn6b4Y8itGZzLcIxuXYR/
ahnfze5TVf9oAsIudLGQPxafwxnxA+ct93lnsBIV+hZ7HgKV/N5khkfB57TUDU4P
d94WYpxSYWjbbZxQqFCiooX/cEe1h4/dpokY7NzZNFH9LI2AQJvzVMYSYGY8Y8vi
anzvdLHa/jmtfin1aVEGWWZk85w1eh1ReNAegPWnCJCWhQLwpOvgs+8QxO8Zc0eW
yGlC1RTh1jrr+aSpuJknityFYkK1Q8lJSvt2ZQ44WQUYz80VhnZWhrDaofdbE+WR
1zMh1XbyGRw2T7S3ekARTjyjppTRs3VtA2qfH2QAw3yQRTJjkYOJJVwbt21vht9f
+5+5y8VPGi1hFi1eydHq4ejkMWv6RXZ3DaM08cBQv/lDLNm2GoRMnP57r8cgC0Tv
fVIdyR2SH5WEyl0SS1QTbnMf7WCALlNDiBawrEa24kTDXV5rtb6SSm1bYcrY/WQE
3GY9im8h4Jl620pVmOwB7vZ8Y6ev3Yg8atc3Iv9R63GBg0+UHeO5gY5SzM9Ob+o7
1JCakIkFVwj1OF7q2gqXhqQFHzlVHsTMp9VyxW0h7d4qW+bwvh9ZxxhwY7mjQTUY
QzT6EHuAR4S6Q7EapKp1VfOBhAsGn70ELmXr+vOKQnxM6sGOt/9ovkhQFMfml2Ft
b+/J93Ymd4XopK9cSrNNTnKTT+1OtLnFUom5UCS1fit3nrEjmNZtGadL/zcT+hrK
eGf8T0WA7OajUhU2zqtC0ueJ8O5ULmueAEa7oDOKSH877bRGspPyZ4tjSZaRNUSs
yNqifbIU6d2XjaPsqSbk2giuHj4GrmUpF/6hMxrbD2MsALB6Kyvz2Toyru2qShHL
DVJlXEs3ivkkgI5hmP9js4suCZ/OwucnqL+iue0dUNiIyUPQvfV0eUyNC5a0nc/A
NpJ8rvFLQGhL/YcyrBIVCdd6zOSvlaWsMLZFghqf+rwre5TJmXGLKjosMFT0vDq7
hzEUuEJgLN9xE6MiPOJlUqASwJasYgsHu15hc0PfqQ/T5WI1KYTQK4aI/JlXRofY
9aMLATRXnh38r+leLZToKlUaBvpl2YUEqQ0amqHoMk4g/FYoDZs35dq3CYUk3QkB
yFtQE8JnwIvsOHTkaHJgxrYUVP6bLLgtsIIn5nD2GVvaPPQDfrREpBJzy0VshILU
qePxnJVEatpMsjnXk6Q44CsniF/qqZirsUKUtUCNVtYfzc+tXunWTMNdKxvnU3h1
y9VaGt5D1rneA2/XBvuXvv5+uqbZcXVvsQGKViBfB7xSWYxrWMGEOlFvU3davGxo
0a63poD1DrvAFGywSlv4nozbWFYru8WfoS9SDeX00D17/BG9Xy0oqbhHPUQx0NvD
EdYx9PBRgCzk5OrrL2Th2U5m7BdPtRwySuwhGZoc0TDin3YXWecelTbFCIEsI2Tp
W9EUnsvcI6gOiSUxAD4eK0E2D72N2A4V5xUdmpiOTs5StEwnCB4muvxsEgv2DFkm
2jj/eqjjY+wWN5QPPIwnRgFzifT3O6E9UlsF4UZzAaoyokFBWKrgRPFjCym7IXAZ
B2t7ZBCedbFnkUhJKrirfGfs5aCYGfCQJcHpFskbuVXGERnDC6bijxJItsTQr3qF
JIbpq0lcXhw6y9OY4+CT2Jwi55JEkugpljK3KiXaIA+VKtSEQ9wbHvzTJUOLydtO
FLYOQchYJ/MIPh4yFBkgMWZoYkf/V/oAlQeCgLffSfinD0I8VbxqB/aA6gNJOiqP
OwDo+0Lfd8pdM0A5xW3/TuQJ/opBAV8nVWVHBX+HQl5jkQUONtepvYZSRninAtE3
EnILWuWxGzlKMkLfJ8fYvZGZ6/eKqqt7YuE01joKjAFlh8Z0I4Ac+VPfz+wJ4Rfy
wMkEnP7Hf35qgB01rHMNl46fcIBT58ku8iAh7lA2L4v8D1HEdNC4uXFAhgpiPXYI
YjXhG141G6LPSJ1ndasBw6G3wpektbUGZLAkR3GX/QUM4vF/Cu1HC3mnzMU1vT6C
ZLy5EqyuZFixFPHMLqnmpzpXkLCm7EsXLwjq1H4OS7DtcoPHoTTvMEwpjQktdV8d
D7Ze4G8XHEs7ZwqaOhqlv8QJugqDcunJcnYLEYfmuZIatzuuCa29NDmJ8lRUOdC2
Cq/lSGdYL1LuXgJNqg6jpU53rcphzwLzsP/SBqFrVJh0MtST8XbCca/91qhi3NPI
sbmJRA8J3at3BhOBRcE4C3npSA6bKqwIvzpk9cZuHpx8YlPXuXlG4rt7p8lKP3ip
Miwu1lQEqUt2yGv6u7NqBphyYZU5OBhDMqlHWGjb09SW3DYfNRg4d/DiRQ9LVids
eDNYKey5/tHtq0FjweicD8DjJdFcxtfVHm++2X9oTMIrnffPCpEFDhgcQWyvpXaX
Nqp+bU3fYBrKiB/U4sootk6edY8MGa69VHOEtTsenyXNqD1x12Ala5tPvusq2U6k
LHwhYqgFIYhLAJM/npze5wgBCmSowvJcarqEUcX5dpsYIWEYSqATUH7OauFc7CFP
q18MnxX6sTsODISqrbFL+ecWqyfmURq84+uK6ltiG2kbMby5t1GeyxFNDTWqmhxw
ZvVKVq+XUrsRsX0/6V9ixfPrLcq4zcz1IW9ByGVMIJyXsHl5jHqW0rcAV8cmhJLQ
srGIv8qoXq1I7EJ0FZTV82v7LytrCpZP3qQkBIflQISNUhl60CADwBruEeXNo+3a
5dwIySsyjUzPRdqA/vCLA9bepUO6KhuTAjnOHSVQF+mKRnu/TSH4A/UR5p3zCeSf
3RfQiNpnbqVdr6U5E4on6aTSBOR5NneyK0x09Q+uwaqXNgjtIi9AsKkkKS45qIQv
amp4I7My1kbRDX6impzUXnQwY6z7MI8Gp8bV7HGOPZ51yVLpbuZolWxk60ebpMht
qBr6LzfWm7h02/F6E1F/66rErAZTUJDyFzkN0+l5swshd/JKiG9Y/1lpjO7CE8je
GYagu9DHfoQjcdsr/NjTgrejk50/WJdkG6JOOZanQ+q4yOx6AudFZYDPaoVRKVCs
AYrLdyy+6ZIUm1hsU+wriFMeb2+6jCjTzuIsErgBsv8LHyrbxLbrQ9B+fL5ImBeX
BB43OlR0p9cLYMN4/C0ta+IZaWuedHRwXpttYyO2Yi0IDQj5erpHj9FNMVQ5i5It
ltd9QEWqP6hXRiDaOOS+UAayYxl0O9Ln9u0LJBUCg0FdyEfCk4V6FHIoIKrDPBAN
KD2P4I7mdQwbSKO3UubWQlZNTCjSizgReFnB2b+mVAi1yKhf1ztQLJeT6j3KRQY6
hZ5s3B9u8llsQwhAHCSpH7lycZqbwNzMvFe14UwH2xdq93hppMfW8ngu7+gSrj9O
As56yi/7o3Ra9U99IYy1PRW3RdeU5ZljERCAwWFbITvH2lkBlJZfPASWf5mZTGtE
eZUyqtgRCSaFD7peGfwhZyq5cn/rNLpBYdEqvJqWXlYjQnZ0VC+bNPQ4v6T6FXgn
QrOniQ0NN7DH2D5U9dKIsqJUI5XBjg/kuP4n8tGdKKm9OvqPQosP/bvVDE3PN0I2
SeFeFGZf7Pahs6VAGcyWpg3WI+1/LSb09DTItaR+Z9NkODKuw3i1uQSZ0oa3gMtd
kh8H6oTQT0vNBe1ydZpjb//jmWBH/r8tmLBkwkzSVvKayqC/IysPPwimGAXoqgcc
98Oe5foipzjhu3AHUxtA1esPEFBoFLw0DwIwo7Bk8xefS0plf4PMc/TwG+79q5CO
4vsxQuGXY7CJ4KFo0mNVMPKFg8OkTOC6fKPzrSqAxLt2f0rtNMSSMFznYjbeMpxw
+9SqCaHAWNBEcIA0SIdcIqsK12sWxF+/D8EzrwGKS7jWl/NTcabY9pc9CWlDPvIV
JNLIVBf1o4MwYzSYFhPyfwwWj1cd+tg1twRI/xN8VhzRUf/jZ9MzfSKQxg7i0Xok
DZaqTCJg+N7CGFlp91gYu5UVmfo5fj/Boil2sbj++A6GLkGr60xfQ8IUR0PsACM5
nCfhiO/pKvQdkftQZ6EWEJ1ZE5UxTYZtsAXHlUfwY8jTdYHBrx/o8bhfcMDYHyaq
KgdiLafUrxpJZhFC9W79za1QMeezsgteeiQMklmf/gRKjYwKQ2lgXDf9MorkkE16
1wxLfNS3nCWRWr3EVEFCBVNJKndLiKGecPJFCbgUGn0huLQXjjnFBA662Xi8J7Yb
y3nFJXpddkO/cfZHLcqXPdK3r40ooF3kt/6BtWJXv7BzmOB8FfEKrKhno9EXcraW
+1ZYHgtFYNpVVj2cr9Wh64pyQTwk9zUEFz15sbcrvUWWKVs8HZGHnEjds2CUJflW
TOj3toPO3e4zEUDAp3vRLqABwJdAXywb5fMtcTwuHaoA3oI2TsV6cwJx+VN5PSZN
MLIhne4KeA57gnX6QGoqtjJ9xOvLE9tew+DoySekXDanSCKqh3VigBMv5MA930Qx
KXTETcV+tXOLR+FtlkK7RErFHHjN+uxbsAD0fDUvhf+peugs7d5p9Ez7YiBxJjHz
p2kf+qna/nMwk+ADteEmexArq66NjjeG9euFutaUUH8FSCBjC6ElJjOr7NTpvW7K
kWRqYaod5xWeelT2jhMvmEEJIdletGaHrFwy49VA+0YFKjTvkvx/NfM0NgR4Pkc6
qDK4fv0aGKpEjl00DFymR+kL0J/0YE2ZbMoGXyPRKAJ3SrN3hUc951t2VMxaaR3f
el4CvyeCe5x69dCg3M2tQuhXAbsyprZy9AYleM0muR1qm1iwjgC5v/QYZHuF+f1E
+E47cJ+QI7SVpvCuQ8YmaHVuSyQuuz0dy2SPaGPJWSTBSE+rHmO+Z/QB3hfCTZFd
GMjsZXlW1CzMjpeFosESxifXyi6PXS5u7KvNHnzXvfYlhUsDhTwnd64il0fbkFxg
/vlTIRjqmEt/SKyjOHnbEi+yaH2Mim+3X1m1NB1hkEUP8J5ttVEsSxtmdlxTTezn
A01W+iyaagBVdBWX/MmGiARZPdeyiC4L94ePKf2IwmM0oD19uigCIDKPCg/ZEs0m
dasVNjouBTHoinshuHDGG769sJvHwMOyJTzPCxPnUR3z2W9eelMUcoXFaxUe3qkL
LLBMMw0mJYJsYn0jPZygm5k02zdPcmiD/mnhCXeDEd1hXapda3cYWrbVYuKgW2e3
MWO7nF6F3e6+i7uc4HxVdqZtSGI4oMH9mUDMc7/TFxQB+2NbvUiA8/oeLZsI0vV/
0AyYSy+dyMpKRkXkjUyjfEJRlyxuwL+ECePQ1y8bpm6e2n8X/ih876VnVLg6spbD
70SK9yJmODncnTS8Su+Gdg0DMfIaxoeiZiVeXr9V01czHngVgL4lwUfLpvewevLy
Z4rmNeSWInSbjaSxdym29e2a0YreJ5sKRaP0HfDw1ZaO0QUUDOXpAXd4762+2kNw
uJ2Gi5wiKTFWbaifqIp9wqZ3PpGW55zgPhYxHGJE6eHVI8SzRBBox9hzwEfxLAfR
Ctur5UXmnETIAXgV0Bi6RcLvp2xv8sXTBbCGfbDz0CSp6Z/qkHW3KN/haCg6YT+/
23VpEyV8NHJ1EsVQeK9NzNA3LJi3ywOw19a9YAy/KDEyTT+QAZB55Lr2mwiRIfZu
OkgveJ5wu+bSe5V5ESzxX6/VjPmbOKVSvNxsNQV70Vt4Ji1TssoELRRG89ajcqRC
sgFxiThSDQg2A+CssBc7jV/ywxjvvYmR2hvJhSYo0LMbah9Lt6yS1vNXVY5sjrGY
VozkC5kQ4dGkH5Oi63sVKu1O8R+XA0y6MPnUYFv0Y/UjWEMjhUvhMKAiRn/4ALNZ
BncHbSHE4a14DJevIj1/8uDAwKj5dv6oIDpwR9g/Jy3Heg/kVod/w6BTjd5zJBw9
GuOgEzG2IVg316/d3Fep996gFxKmC3TvFp1RfkLoHzSfnX77ml03Wy9MqMQPL8ld
9fsl0jhu5CgG3YfeDOAC/DarzuJgMME9ei7i040ooP8xjdkQaDKAq7l8aS/k+RBC
iTNgjxSsvIUTKvmI2yNeNJHfwAFq8q6pQB8MkVdASlZj7/pSe7Mf7uUHd0W0Y8YQ
JqPpS6/lsucfZWp71vCN+NWP2kU9dhUZSPbAaoPdWSJRzcD6kyt9Kw2SAy5vbcTi
8FVEO7NTpHbA+zIhjfY2Kf4GdIODPiWKbw+OsHRc5R9UzebGQmKFLxpH0AQPSGsT
xF07ZAtRhtq19BqVjCy8QRbNuG7cZ/XBGAy+Tey80co1pD84laRG1YoimyPSxl2X
TIXkvGOHYFOYLBJ8pxOYTRpesCNN3pKqDZVBJzIvGGprKulJKVAYPsQ/cbpzVLJf
yQgWC2VTF/wRpb9HfjH0sXFZStLWmXcNUs/QrRdSmlPlI3YEGcrqTYWiX9CuG++f
tL2qbwGRCU2PSQsrrmb8gFzRtCw7a8Cdtkqhnht9aGMddfQ9ZE5pfDOkshln3yTD
pfwCsjbGs6DqRzccNNLMQrgxJgKNcjbeESZJB/vnzYoVImX2zXYRV0dRlZQOkwtU
iGJm2IRMfbL4X1BYgWpBcwzucuJwpb0oTPTNV1HEFTup2OfjnXWdNz+O010kkqIf
OgGXpr3GRNzpe3mQTvnaPPs7v9WB7fMa4iNRiCoDvkC5/anOcc4sGQlXsyiIsiTC
L4ZGUUBgf+7hRIW7ZuSYMJ2ppwEzED2mNimnkLemJ+aYgRM0eIJeFsQJMbYRl27y
sxX4cYkd1GDj7Z0cWH2Tizp0Ku8tXXFpOP7fkhmLKsLG7rnYu90RkMzmFfz6Icb7
JHj0qPAy7nIeBT8T//zr4dT4BFQNWkKOd4oGFqt+X19ihph9XHbzx4KOawmxhNU7
7MgVYpvpg37MDSir3LSE1FuPcFbwPKb6CD9guLfKqznQm2SyABqtv69FTNQZviQt
7ggTn+EBzvxjjoLCUpj/qoE/MqdYreAQsc/5Onc1lCiN+Med/ASEgdYuONcnA0Ek
Dw7r9kcThqO4nFVJosuFennHJA/wIlHGGZiqskROW+bG4kRiLBIQ9T8C62mchY8G
IJ2WRHHxOt4Gnxzsh5m1Cn5zDfcwoZRqghUI6W2lTSwfaHxxWGYGHVCArBpTRZEh
r3+8P84TleY/B9MY2Z0HLvyEJNqfH3wJm9JuIg22EcKfZwzwf8mh0eBOWUJK1VD7
IetHjWOqyQKpqGbAhWa0jwoO1q1K9ZXyT/C5WUu1P9OOlo8vLT0p786+prktq4XN
CSgwZDAOeb7thuC5Qq5rQ5kZB4DMt+J/9pM16rOJoGeTvpypWn88hzZtIQ4ywfn4
2MKYQrIKJu/cxSWS/aVwNi3aMU4p40So5DMxORPmmHBiRa2ywgYve+6g5XPDa4Y8
sO1zgINH8iQT7VMvQ2PlAStebaycSBIwWmxe4+ZYHd5Y9vt34RljlV8b0iMVZygW
D158SIviM1erF06G6GhjbB27SadWXq9Fb9B2Qk8DMqQvIcLVNi5H2mm73Aepz2wv
DPyNBQsf0ljT+wc7AN818z50XEQSX4zd5gLzW5xEFHJX6+raKBtOZupCYclhUrkr
YQraizcSQcM4YNKtcQvy+O8QTRuojmuKjuhqjk/H476IgyrkI+Yu8J5mhw4l69XW
UGs2YSHm8kp9Y0MU+yEdZPz1mz0zm6dkjFT0RLiGa8uoB0D4Kh0RUkwbtb1U+pVp
suBzcMBiAdgu/cti/qvfkL0tEXxduXiiFQZ04E0CfF5UOuXqzygH0Nel+maI7ctJ
5qWnw4ZuWNHHaGkd/RlTX9GlJ1Ds5B00VGw4ferT63/uh3FRaYdLzyh6N04yQyGZ
9HoF2sZMhZuYhbzUBpbsgXXX0vwhu5mbgux8EYaYKw64XEAs6HAFVvwZz9AAKDFO
9FNUOvc5/vS4b3AnDc4wz+yOSAHo/Wz42bf2dYs9SyfiHJbDKpEO63E08Th0szpv
8L2pzMITB+Rp1jvtBNKNlfmKAwCS27jHE/9P8VIa7xtiYmfH6/MxaCZO5qxqkQJI
xo3f1nA3NIMtp9+lKu+sKKiop6qqlQJR7LZfd9t5wZr6JdKvgVXXwjULf3rp+uxF
4WbnsQVojbvvFxQcDdIzuGH/7lqLKuLbG3GyrGXdhDmUbUx6L9aPz/5ctvqEa6pB
esJfqC/bfELqmpuYPIriAKAnVgimpTGJCcm0+pufbFcRZQT3budBUnEqtpfjCyCs
R4uO8DYJBEv+o5+tllk6ZF1C0MBRU2x48VJZ+4YXowrpVhBIHbMcgio6vNNM0EBM
KuHUT4GH0sqEEdgXtdr7PH2goFupeSomQC4uN47jYRwemWQE0fdMnTqDCQRjr/63
NM8X1uW3Mm/tot0SjkCpYpMpGgXKaVjqLE9YKe1sJNl92Yzb+yl5XvYbxSQRRTKr
b2gJrWYjfw/N6P88CLxtFbUdtXrpvObU449jpNDduEJfPmdDINiBJkpZ/Ldo8Woi
K2vL7Bz573BV0LxXTzRun2nvcmpq27Je4kyg7X2hNk53NrASdwwrprtJdNzGxeoF
uxnVYxA/fl//9d0jq6wStWXI5OiOl6Wg2bFu+QVYBAXYBsmqL8Y8B9I4L7Z6muRj
OfFimShjM2vKZKg/xDwIHANG6QWYWxhlJWNJx9L4zfh5llR7gPdz3Lg4791XqhLt
9/LG5jAvn8snTH9hlMnAdsdUzZSzhim9QaCVp4/Rr8WeOEKoAAFXDbsIEa2/jU5c
988++OdXdJWoJtXgu/Rh3k+tm8bIO+m3d8GygViethBnn3eRXiSrH+L0Q4Eqv1BS
lBOqyuV6bmEXsxCJ1or5XFyZsYPAaWwpXM8SCDvDImp1Jeu0P92FlZCXbLIXrKDl
6+X3AanG0gigAwNKO9aO+1YwfbH1uLn4mIOBC1mPWuzqYjDbFKtpsETY4F4b2yD/
l4KGE5ad/Nfo5nXQsRqLBmukYNmqIx4chZLIdN2+RWpL14iX0EmBE0+5eS9RJixn
kgZxaHgoj4u47sIiWM817kCr9SOpzI9Bum2ON9kcBs9608nanflxXCgTZyExdoik
XMXha6zLYKOEITAkm2jG9l22XqLN+572Fa/O/riKITZrav20RU3KwzsGRN8RxFwG
/kmIBKgx03HbhKWLuVGmCzkmtWa/E89txrpocbL34lYwoPOPSBbet8kmm9ivRtKm
OnWbyP0UjvS9JExHiuzm+KPWCXuFVhWAYyxkgHywRgGdD2adN0HLEvqgKQsp7mfM
4d+2XUF8C+rrj+GU8NnBPEgzpTTuJ+3SWCuTYJi6qTcRDa5G5HO10GfbdQ6TqvH0
F7Pd+l5ukKV/fuKQRynaDFbLu3/KTeOs6MkFCAEpvNk7kYz9Kjxnv9TYpm1v6da3
PIqISK/5NajI7QkgmEnKXDFauA5gkddJQVAmYqJbWq7oBRYREGQCg36/Lh1Uicch
gnIjGEx1DlO3mVQDEaWK0LUXdPAyPlhXeryk2TAk3pTahFM3/ZlZXveYtHOY03Xq
LHXO7jnbQNwEkiqnFJSDaIwW8gUOrHskJfeUS5eMQc1D0E2hR/zlLVG1fBSURfGP
jTipk1MwIPHrR1DVzIsLysn1n36c2oV861h2EUjRrEpvVCcHKnrrN7/wfzeMEeiY
oA4nkpCTLrRNOr+Jx6+smPzCNSkKu7Xwf38ebd5QjrPb+w5PtQkmtAZWwrrGdFg9
3QM7i3IY7HenoT7Pu1Vbc00ecNNOdUfpG+UTts82kWINxYAbaT7Zvf/kKMziexWc
jD5NuWx9IQ8CC/b5WT72UrieuiBzMe27JtFmOk0+Xws2vBFNjeiuN3ESlO1V7Wwi
TFKHPT5w4dB+gb26Xr0hwxilhhG1WaKfGiiFIJ7PAwh212tdkTFhO54bQCBHcnMl
6/BPdc0W4R1/SZhgMVm3JtO3khxltvj7cFmp2GUgj8HV465A5k66PHKQShzYFYgX
2XokwWMkL+817eQRcnEHXSjwY78WhOn5+VRS4JscokIKVj5v0zW1tsQYmhROEbJ0
SqksCZeYSj6O8DuvcUkavDdLokVIwcNVidEkkWJ6Jrkvy06KV2JErmxzcdo5Vn2C
C+39y1XZYZ/kjK6xC57hIvmtY0EcJdCpb0sssW4sPOuR/i95hLVMW4kQmVdjRuNA
qwwSoHNPOacwDJDOwNZ3NCzxdpJXzXpKPUGDu2T79/wAJSz+rKB89/JqR4Coh7J/
MicoHCUWptgw9pfyanibXmTQgmnQjZYbi6KoEdTOFyZ5SJ/ajj6HFjr+Yc/ZvQk7
FwMG58LeSCejp69EruzFeDDxSWTB+yk/R1NxikyQ6J5yqQb3zdhbY7Uu2gwe9e6e
TiIU/ogFLbS3eUQMeDdU0OS0Hmu+4N7pKiHb9hArlrulmv2iwKeUlRopuZ1Oqjkf
rAW7Qv5dWBRaDVr03WC5n2CyZtmdI3qA89M8YM319wPUbJwmXVZGi2uFRDgoghxf
SHq/Y61bCilA6Ut6zNN/6rGFck11Xn79CG/per/EQ0ZwfKHiLhXgipxHZmztkzQT
WWFgm3+l5l+EcCSStp+WBfeEHraeAKw5IucSCLzjJyVuTUCTPLnpM0WLZX8RnxWw
21CjqAMnr2vOqYFu+OEMA/DcIqSqYI9wuujzCKjOJoivKXofPjQ9GFUdi55Hq4BU
Qza+1ThAA7wFBhqQ4egpncRB7aEmb30u23IXcbkb8A03jAXOUUXef2Xj/aKn/ljj
3T+L+esinL1GX/U5Nq4nmX/MPg6OsiIGjnVjaVI9jpCFelKXxq1DsIzxh0XWcpPt
LZaC6VjHtku5dWIUebfzuKkiK3sK9z7Uk3bMfP/9vJlyXtsS5nC02VK75qm1MlB6
PKex6DSHwR5XeyDUdKCG0D2pqlbbXnTAbEU5mY0aFuVVwVrjM12RSNgAkuM0805i
TNpiZM74ruXpLr51uGCVBt1cpLeYBaJ6QElcmA9wQLpVatbSDf0wV73AGHdn7QIu
JS+wLdnDTlYGjjrVp9NaHHrTO/P1uUEIszs/c1qQY/GVslEkv2GOgvApbZpUtfCw
OrsQUqxNttUfpEt9U30Bnno0KKVDk0LoFOyRS0LnbzoCEHPkibzKOdPmwZQ1AKFf
oXla2P4GHRy0SB9xhRifyQKcjqT3qiAxSiTuZ8X1ta7DAPEepO2UhuqcqMgavaY8
RJIFzurAgkgwC5PmMCize+FI7fBsmT9CGAedFj+jPrQmFknLqyQcriQABWZ/qZxx
Eh3SCoMhFYgzHa8pie3gkEnKcxoeuwYJWoW+PepZgv7u1+NInCTF+mYbyKtEWl6M
dhzXQCTxkWQbtkdlDix2+d4gNLT3IkCWlvlG+hHdl+8nrZU1TL587pMXHQByOtiP
imsYKHgWPyQLrIf1CSYnNP9CL2Zwt9qjMxyRhoSz/kpJd9jEZ83T0Qw++Gzv46u5
UUXJIqAg+6ctncANuoUu+vry8QpNqg14DoagfT3IxthYY3BQDMOOTHrRQhupC8jO
gks2z3/txBma4qOubptluu8wb3eaCBxNHhHU8q3ovPQICEO3kODzIx1rVLGslMLD
1dEgYdBT+POkDp7RIVc3bOTa0uQCb72YUTOMHn09QlN5+L4aNwG+ZCRsuzLJZUKG
RJ46WmIiibu7cYoQMNF7V/vKcQbOzjRFJ2H+m6TptI2M+4vxH5u/XjTzj29IH03+
Ma1BboXMsB7oYHJKEl4o7sLd6hryc1ZcRSc3gws9/xgKzkGCgrhyte0wCy/fDDLT
czmg/ClSGAXkKo1MXxUc7YzU6r59qgv+ZljKaS/cxGFUR6kkWV8dNZNvNpM4Grbk
rfy8xXkBs/xgZ6cjzViWVbT/2ezbfX0tE1scLJmQEtquKGyEqZTlhrVHRhlBwHaE
FMkpv04s5rPJaxYlgVUc/XcM3/6J6Yqo+4v6IQ4+8QcKc1psu3s+aFcVzCO9mo2N
S9CZwqz9QNQvdr0fVzYTV6ts0nclaeFreBZ7FdXh6xmAX5mE0m2e+mCoRsSUKNQY
kdRyugPDO29pQF9kyqGM+iw37UC9IgKnb51ebZGXLIo+4V6qeccj0nF29TbZIqzN
M6ujYJbyLyAsAj5RjPml1E7PS0I6dhCv0WBN2Ert0GWGwHfKXWIOHYtBkPox8eV3
yUfIL91ld0OU/vKg4CTlVXrN8A74yD1yrwG7yfKeq/VgWSnoyJOAhMy+FylQ8O1z
RJwyYhj6Rp6fA4jIxxAIjbsXowjKZl+lYTI3AG9es59jMmVPFcJGUyWV+siCnCsb
bddpuZW4FG4iTOyOtDplFZOY/hW51w5zUMV5hLw4Z/TJj0sYGkxyfJPsyfL327H8
2vajhiqsPWFdVN+EEdoTPoCzPFXTY2oVhjB49l4+5aRpzCny3fRES5bF2EvKbqZ2
gyANk6wloespjEM5EFo+AGOE0hxQkHJzPBCK/EDfgrf95AW56yt8lSMRPnSrPcFn
LFeRhag8FzJbpgMKEN52LfGngLV4KLeRtCRUodseyA4LqOSynyVQIWqU5jao8EY0
YVitq41VxRatzsmGa/raTnnwgccXo83NW3439uSufPfR+wEJ6dObCx0ikoz3FHA2
9NtrC1h0euY4F7QhhHeWJxfLsGn12yUWyuQb2N9oqFVc6RFf0LCBtFsoU7D1PqVS
/ELVfmPNcrGvaTz+W1DdlOZqmUKMDPQLWfdoYYY0uZQxbKoguKOsCw/rWp+RzjOH
5Tqp5qzObgeduJDOFie1xBuFBVXp5hP2mWlcOu+4/XI/R0AiVuWn9YqY7ycU7QhI
cEMHY8rdrzQLXq+AdICJVWIJSxuLC9g2fGVZU7682l0wpnLrVfy0DMs+CdF/jOmF
+RsCm8fJNcSmY1FKnu4jxFKh/KlAIX5nytPnz/pI2REj/iq9q99JGbwqtwKaHdzA
X1inYjkD//AiuaTsKkeAAlx8vSF7DwUDrCRTU2V3YyM3/DzJRqPUQ7tURsXhiuUZ
gqPvp/NLJOfM9KJvKiIoymQYyaiYGnt6QZSoYhZOo7AYAZcuSdpmDMUWIvr/uUEH
33Yu/Ghau1Df/lWBoaQ/1G8F2Z16s7DOfR832d4AMCcTGYqIpfRh4duY/IiVwvdp
Afh+z0THHY1cfpSvsDLhMzYtHdmBi0cuYQgWWUs/eRzSuSvUtWVlcrS/N7d6clU2
ks3A6aiKQl553o33rqiATlOhfXbKYlacIATNOuMhZMJ13vwbISkkRswCUeYBevRS
jccm5jPsqUYcBYEqQcJzZjwvQv0CXy/m7WVaKIsAqax3q4EfsXf5NxMevbL7T8IV
8ylLUUKwyTqtinE4RiL4BE65jeQO3f1sF98RhckPB/cQwpsEL+C8MndeAglmsJMr
zbOHGql3uvwYnM0jZ4KCnL4nkPRa9G1AeoBaD8CN6CK1SLRbDry3z021ZooQnpY0
zM08InEhUXSpfh9847PJ/TQNgtvvyUSM7Fr+bfvY4ihVzhY6pujA7hrtvq3Lq7B9
0pt4NWnU/lBp0Kso6Z9DD3p8qX1uOFbF9YEChESVh/gPndW3FQKK88uSANNKNxn+
dMw+bm8ssNvXYgkqSutznY4bkY10QLz8NyS2ROJTaG+vewADejvbeTIELFfQT86r
yhZVjy1L5CLJQlrl9DTkPDassenr4sSfkgDiIL0rpo6yYvqSrclGcnvro0oITXpW
jHChTMzbb8vDqb/HQ/C8Tx1f2YOT8UdnpUP2PYcKsj/NXU5LExSVjLY8aJuLfLWk
HgaVRSqZ1MdWiqGmzSqjnZOJ4wQyPyBh0wLeteEDZQ3nMd3Xf+/QNBbBtyMgUiYZ
GMQMzIx2+jZBXjfOti47LZ4d8DmQve3Q61+/pE19Y0TO41Dz+gQ/BYTUMPiuAenc
XiwhXqHW6aOF0gepxzsM5h/BHse6XVEh9yzIhhdjHDRdjY/TGClCkr5Vf+DnTUUF
JDs5+k7dRL+HLmWKs+j0J8++e8kqvf2UVi4V0/2KgD9cCU92zxLzClhN0uoy5eDU
16m15++WRuTOhF3Y2N0Ftt6TaTBJXI+BkSvQ0cbAY6hMvYS8+2ah67topC0ErAWN
CfWp0Fj00rZ6VexxgvkbccK7YVjJKn4lCRFBybgWqeKaqRG60CPW957kLQYNzcr8
2JzsBJnC2EdDZwWfJDREW3oFLjuirovMkS1Z8gbah9zCMNrNHFZkExBEhFtJ5MpV
BRFO3x43iyxCsfK7t5QGjPDu1ZKtK8IHXZxyYpc3H2S3H8yefF1DfCDFMra+LMc1
64EpO4YMOCmzwkElOaVSnDR+UOTEOLDqz0OjdA4QQ6isBXnlfQRTPA7aJyjnzqmx
ZXsosKc9Ss6FYUtPmemG3JETFtI4R4zMTspCapir3pZUJedFRMtszvznF3CVRQKX
MhnHIJX4Jv1GFS6zJuUdryCJX5gyWPSOM0iX3dvtTglka9FewCHiG8nLIJAASSHX
VKb/LKyxdDWO3azpjXre9lo49UZhTiBnrM7sjCEO1HSoAByDXgDvs2K1Kj+1wPJY
Z3fY6el9DZjPgr4rJ9Uuji1+pRTIbe57SFKeywWD42C5qxWCeSyVUDmTSUr6gGO0
/Jbk7wQkJGjfaWsty2c7BiNJCX8QZd/99Xmn1zbm9ErhVKjp8hRjiZqCdt9UR105
LGwuuSqIQZSGQejpMRYHTEwTejjjJgoE28JaX7eQlbfGARsBbBt37toIEaF1FQ1P
L47/VDc1X5JADmWJaEcxv924aZLod+YqeVHGDFRSppkuM5Sz+S6dEm7hJSTFLo2N
r04pHGJA2FFAv/Ri2CLw/pVT8oOff1wWWdHIec7dGTPulo39XPy7Bda4N81L0hVK
dJj73mmMrqW5u4eZka4EeHzZ/Dia4rllRjnWLLhZSJbNWeUZwwFa1eBzKrUGu0AL
7bgCtpDwetXVbCipK8nZIfYmZfpc6gRk50FxN8+pnDmQIf84cBrMyTRl/DDdiQZn
cbaqlGeDOFVpSe3xgWYXhIqlX62q9ymOq7KhFffFTWkPJWuSdxdjfBD4/qdwPd25
0OjtRyrUMwBOZJb/yjOndJlb/AdNxOYOOLC0LnNlp333axVdnDgMFvasGX92zdOm
Nefl1J5TDjO31U9f93Id8lfQT6dff4mZUCINoU4gdgfX2Re+LSN7afZXVD5JTilD
Bj3YA2CYhJzmCSdPkus2tI6aYrQSy6MGjfJmtRzuoY/Q4p1NRlnv5Idycp24fQlx
aGso8eN1s+2uG8wQLffvFUQclqkejD7PpP37f+j2N0+H0CK7+y14UONv+hJ+6VfN
Ygh5cFDgMWEIhBQ2uxaGUiXw4miYw4+EGCLRpeepz64oN3USyhMQSu2pISy7Do8o
xuoRaT5/W39s9klG/YbS7efv0NGYIh6MyWTgc/MF3jxFDZ5KQprRh9ALHIqHzhOb
YQeLClSIVGvH2tUTgb5RZx7X8fd2R2qI3E7eRc9O+xPhXT1MQbRAa2m3aKpneNFn
n8OSpKTEzBnjltWLKOlijPQbqb281vwrfcWoJG79mr/pDjKpqADFWcklfHt+bmE+
3PcRRQzdCoYfH7FMbcqUOLqImXp4qb4hUoperxmVj7oW1xrW7ZamGZiLKEGxlrTf
Kaz4kgL0OH/WiisYzhbEDBZJWF0j6iU7AdtVG30/9jwg3hTqcxLaUQmn5UcxqFKc
O1HsCetYljcZD73CcI5/3drEn5BY3hyd0YyelXfcviAwWK9xpw2suLzjyOHc9eAD
10MS0bK7k4AWJYrWeGPH2iw/RYBt26jTyyYa7+h1oq+ZXu26hz7ocxSe/4zAOKao
IlKoIoB94pqshp3sxgXK966FF+aNAjTckfVVzq3FBoBVJgk4o1pxrzhY0n7xp2vT
XboxJXIW/N/hRsY2G3GO/zuu7pLJXwGyJIdnv9Uhl4PDCggOf0hH0Cwfwct819lr
fyNQal6rhCCGxm3to3oFTqopA7hq86/fhMa9BevGgNC0Kydiw6+eHU8CFJeYfBQg
YBa++2NNlFy8dM/K5YGF2XwNq04cmBQ6ejkAOxZDRf4wOFLtmwJOOQ6TFob0HA6i
6nP2bAWMyuEwq5A/Qfa6EuzHkhB2JSCAkkShjzHtlhdmgKJKqjkehfcyBJWrMeYd
py9HHhBmZpiFfvYbIJycYeBJtKkjJJg0GkKABGKjj6zWcWbMd4Z23E7mV9fKlpto
Cp1gta3JU8Qnr7Oy71sWdguWkhoBtxcJ2Afyiiw6AMsY/091WaI8SmqN5JYNcqi8
SjYhKtEudQmuuxnsK05GZiWpGqSDlIZ10xYg5i3vqi2ajZrqQgUFltLj0xihFbeW
7RofVSvB2TOASqdALPUKvDcOfo2M5M1BTp089VLt5fORO7iWWIEw/WjK7BwFBAEr
plVpoJyBDfn4nncS2wUzO9nK1cKY84hNT6Uk6Llit1W6lQOZ9i9y4PY30rxc92gL
S1fOkoQHUyBiaVnODTmT2Iwjyi9fIboXvhKWepN0p4BEC3F4nAF2vwd2dR6ut/XL
bim9x4ylJOAsnd4FK1D3qVxrYOrEoXap6Y9WnPyY6YTn3rnuZjRU8i3CG+r9obql
7ZdEGB6rST/KAPupKyKFv+RIms+cs4FAZeTJ5Xc9mzFYnI78CanBIRDLrkg6Iof4
fptX8BcNADu4ScfHeD94Z/VU1tNby4cArNTH8eKRWeJ9IBUWY2Ud+iPee5hNZTSg
UARbTBE+MmnIr896B6pD+NRmWRyMM35GIGoieQ8XWQ9sB7ivJZHs82teIGsclCMI
E9sOdQ1Rc+QxuOu8RfD9PX0+y5FoCwhdQw7VSL9fwbwDWMuhOE44S26Uz471MMFe
LtE57ZcrWQGGRJyh1Tu1uGKk2cQJjMhgMsL1B8YWvZAawwz3cWD+27BFGjz0/GgM
Z7ak7NQwcQJBuzWPU6CsDbbrlVlJGogdonCtRitSU18wdOtoYfC3kU9ykqSqPWPw
PqaEhOYRYGpHpG7cQ5P0BZ9JXAxYhZg678s2PB0jigkLjXYFDorhTjoets3ej6Zi
+e1jqGBecQGKwYjPqb+afVisGxWi7LkrR8S29/WmqMa7kohXo9fa4F0cnxT5EC4r
hNLesS7CZFftvH3K9HhypFzlVY9LXqJZd3Be65BcwEaLIKAAsiBgvfWjKmdW9YYb
h8hT9vl3BXaW3y/9VIrwEuGfySeM1ODQIxqZQgI177wWSpdZ2VHuhQlR40WSIK4S
kStSAcoKriirst466gvcu+p8NgO5XAMVcHPRRaCcgobs2lR95uXNJLD6tr03vJGl
672UK0C0964nf3hODakK7UlG6EXBO1wDEZfHL8RDPfn35TXRXjiZDAoT/3qFyCU1
/GcsKKuBQ3isqa00fahr6S9ifMkClHvNnmz6ZAP8oTilE9PeSeDLPxpE8ZFPcV3L
pSLhbR271YJe+HuUX/3lPY3ZDMW8C8LKnQn9pjMkfLEZwTS6p9JTN0HdAnPEXpfL
0gJtWyJFr4OvVw4FICzIpAHh29soqnkyJDkBdEwv610TKFBvoomEbHQQR+F53TKw
fPgZNxKE8QKVuPuCEJfKiaf9k/VRpxQfbUKdnttNe/M/nOVvArAd1vaIKbnBc//K
at1eegVSuK7fAuLSqApArXjniBKwsqJ/i/2FAEpagZtBok2lWz1SaUEj2QUfhHqD
W+pzeej7mmWNBCVOi449R1C44D/QEjgYFCgQuAadMroMMmnb2R4sGLhRFi0PQDGX
fRvGXn71WDPE7zHO7+7ByP+Y9evJ3poAmTUC2IQ4FAHRu31YSmIeXiGkAS8+yLXw
Qy08a33I3NyZ82m35rsvODg69Lce87t1d8lM3pyzH1IO3wqW8YNSGtl3+3KE4/AK
qz4daEGhdr4+CFsrHKU5dlUegh3uVaC0RzbKSPNnxKrNo3hNZjaQdNbXAhJFndog
D14cQWwreiQzvoMvabGOFN2jrPqm8BmhLhER0oRMswidt6pDH3ECDOheuU+an/D0
Cblo7JRfaBWjEoEqUlWhipu8nDdj8cFQJIIsArBfyWE12X0rrYpWMxKmmIsoZI0s
A77iXmMtwqZnx5PgEEyw6N7esIfGEOf6GNjgGk5a7poQYZYlbgCYNsZHtHV4W6p0
qqZm1vi0xvSoYVLzSCTkLS6xhQaxVq6jSOp70SKC3N6j4X49xK213NBSrvmbXQFl
2UGbocsWYaDLKLz5Mqy81/OVLZLA2TwPDPXsDBLN+C5k/vbuzDrJey6wZHgF4jgw
zAiJ9x20nMjMdIsLJrzLQBO9lQdQk6Ms5ooYBZeS7EnO+jA5hcouKYaAtr4+2FrK
5mB6zLwhBQaxlzzZOVgtdr+PuJvtz4kWKLfCK/q9G8489RfJ5Gg0ehQymHIzF3Ws
moZFsLLKm+vB4Mc/xd/UQSaEASKrAfaUmu770R6fO0gRIIvCnbSCDtJy5RV4iypf
fCVEOYOobfXCEeXpxAMfFpCNLiXB8W0MIrXkJ2dq1VTzmhlNWZTr6JtTPBXTEqfc
wS7Tw8CsLTfs6nGl6ErOGubN0e7vkx53wcUfVjkIeMfH07coq1oZR+sMgVFS0UP+
ZqMcCaWJDqjFk17NuXk47A25xCWWeYhX2vmphUW2eAIn1Gfl5lRiMeRQTC55fJoz
BKwzJypjY5PhjZlANOvc6F29JuMHiLTDjwHQGHtmmTJOmPXP/MHxyMiJ5L86J2x9
ledFZglgeHkp35Ld5e3eAw1Rpq+OB8ZibosyN/2tqtO1IoevA2YIVOI1O9rBFvpj
qVFCAGD+2XX+Sj7w9uGHevxLQqoGz9yDo0rtJ/Y7E5ifbcaoNfn3TxWolifSfO+7
Gro2x/Hj1X0NF4tfcooGwdsUtCixZUtpdpv6g1sU0FNLn0BfFr67DvqZMY7cYhsX
yoZLQ2KfCjUWfXci+s2t5gQ9PVwini7Yh2sRgCk0b99I4RQpVi+LDKv23jkCU+iO
cbOz/V6YtpbwhKcsoGMspSYcsIoVv4CAD8yBmVL01qAkhYKDRjiYD3HBytqhCIHS
A90WSimAUE3yCjMip+AsirW36O1rulAN+qX805bePnY/U4uL8Pcu/ajbHrUOnv2k
VG6blxJzpWlmL5IydDksf8/lWiUF9ZH+SxJAuZfUqV6FPLbEACpgAkIsvwTtRjg/
psnq8jkaG76iPS4AP1ogRzzfq9it7+KCQ0rN0YFLdEUSb3nV492qeB7ga/o6KW4f
afqQGsySC24Uw9c7AfMP/DHIiCov8mXteth/fKsuUGzBGP8Ae6tr+GdTpxwXb2lK
WBcJMotB+nYVrnuUMV6Z+9pw2J/EzPUhWsd73ECmSX4W7+Dlx0nyTSl5fztYFDZS
aFfS1ntXg50RiHMmm7uyazoUbmL0N7IoWKfhER604bSC4AtHdkgOGRYNqRS6rgQW
qJL6gq/uG6zznXR3wiudJ0fdEklIJrsiVB/g+xTi0mNt9iR/5J8q6WN91lwVm2TD
g4WmNw/dY440b6V50FQs11rWIueqkgsP5w0XBy9l3wghiiiaW37Y50ICzQ8rl/xI
40k9Ed2Wxv+2kCSqnYbZXxA8iqHUbwv6uiPGnleSEQ0=
//pragma protect end_data_block
//pragma protect digest_block
AFtU809I9AOZbfu2pyxADfLyNRI=
//pragma protect end_digest_block
//pragma protect end_protected
