D:/GoogleDrive/IC_Lab/Lec12 APRII/CHIP_APR2_iclab134/home/RAID2/COURSE/iclab/iclabta01/umc018/Lef/umc18_6lm.lef