#******
#
# TECH LIB NAME: umc18
# LEF FILE NAME: umc18_6lm_antenna.lef
#
# This LEF is to be used for antenna effect checking in standalone Wroute 5.3,
# since Silicon Ensemble does not yet support these features. The antenna.lef 
# file is to be used as a supplement to the primary LEF used for place & route
# in Silicon Ensemble version 5.3. Antenna effect properties for UMC 0.18um 
# processes were obtained from version 2.1 of the UMC 0.18um Design Rule 
# document.
#
# Document No. G-03-LOGIC18-1.8V/3.3V-1P6M-TLR Rev2.1 10/02/2000
# Calibre Antenna DRC version 2.1-p2 11/03/00
#
# DO NOT USE SILICON ENSEMBLE OR WROUTE AS A SIGN-OFF VALIDATION FLOW FOR
# PROCESS ANTENNA EFFECT VIOLATIONS.  UMC's official DRC command files should
# always be used for sign-off validation of process antenna effect in your
# design.
#
# $Id: umc18_6lm_antenna.lef,v 1.12 2002/03/06 02:13:21 julia Exp $
#
#******                                                               

VERSION 5.4 ;

MANUFACTURINGGRID 0.01 ;

LAYER met1
    Thickness 0.09 ;
    AntennaCumAreaRatio     396 ;
    AntennaCumSideAreaRatio 396 ;
    AntennaCumDiffAreaRatio     PWL ( ( 0 396 ) ( 0.359 396 ) ( 0.36 999999999 ) ( 1 999999999 ) ) ;
    AntennaCumDiffSideAreaRatio PWL ( ( 0 396 ) ( 0.359 396 ) ( 0.36 999999999 ) ( 1 999999999 ) ) ;
END met1

LAYER met2
    Thickness 0.09 ;
    AntennaCumAreaRatio     396 ;
    AntennaCumSideAreaRatio 396 ;
    AntennaCumDiffAreaRatio     PWL ( ( 0 396 ) ( 0.359 396 ) ( 0.36 999999999 ) ( 1 999999999 ) ) ;
    AntennaCumDiffSideAreaRatio PWL ( ( 0 396 ) ( 0.359 396 ) ( 0.36 999999999 ) ( 1 999999999 ) ) ;
END met2

LAYER met3
    Thickness 0.09 ;
    AntennaCumAreaRatio     396 ;
    AntennaCumSideAreaRatio 396 ;
    AntennaCumDiffAreaRatio     PWL ( ( 0 396 ) ( 0.359 396 ) ( 0.36 999999999 ) ( 1 999999999 ) ) ;
    AntennaCumDiffSideAreaRatio PWL ( ( 0 396 ) ( 0.359 396 ) ( 0.36 999999999 ) ( 1 999999999 ) ) ;
END met3

LAYER met4
    Thickness 0.09 ;
    AntennaCumAreaRatio     396 ;
    AntennaCumSideAreaRatio 396 ;
    AntennaCumDiffAreaRatio     PWL ( ( 0 396 ) ( 0.359 396 ) ( 0.36 999999999 ) ( 1 999999999 ) ) ;
    AntennaCumDiffSideAreaRatio PWL ( ( 0 396 ) ( 0.359 396 ) ( 0.36 999999999 ) ( 1 999999999 ) ) ;
END met4

LAYER met5
    Thickness 0.09 ;
    AntennaCumAreaRatio     396 ;
    AntennaCumSideAreaRatio 396 ;
    AntennaCumDiffAreaRatio     PWL ( ( 0 396 ) ( 0.359 396 ) ( 0.36 999999999 ) ( 1 999999999 ) ) ;
    AntennaCumDiffSideAreaRatio PWL ( ( 0 396 ) ( 0.359 396 ) ( 0.36 999999999 ) ( 1 999999999 ) ) ;
END met5

LAYER met6
    Thickness 0.09 ;
    AntennaCumAreaRatio     396 ;
    AntennaCumSideAreaRatio 396 ;
    AntennaCumDiffAreaRatio     PWL ( ( 0 396 ) ( 0.359 396 ) ( 0.36 999999999 ) ( 1 999999999 ) ) ;
    AntennaCumDiffSideAreaRatio PWL ( ( 0 396 ) ( 0.359 396 ) ( 0.36 999999999 ) ( 1 999999999 ) ) ;
END met6

MACRO RFRDX4
    PIN RB
        AntennaGateArea              1.0800 ;
        AntennaPartialMetalArea      2.1610 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4814 LAYER met1 ;
        AntennaDiffArea              0.4544 ;
    END RB
    PIN BRB
        AntennaGateArea              0.4816 ;
        AntennaPartialMetalArea      3.0564 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4526 LAYER met1 ;
        AntennaDiffArea              1.6200 ;
    END BRB
    PIN GND
    END GND
END RFRDX4
MACRO RFRDX2
    PIN RB
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      1.7924 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1610 LAYER met1 ;
        AntennaDiffArea              0.4544 ;
    END RB
    PIN BRB
        AntennaGateArea              0.4816 ;
        AntennaPartialMetalArea      2.8412 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4922 LAYER met1 ;
        AntennaDiffArea              1.4700 ;
    END BRB
    PIN GND
    END GND
END RFRDX2
MACRO RFRDX1
    PIN RB
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      1.8572 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2258 LAYER met1 ;
        AntennaDiffArea              0.4544 ;
    END RB
    PIN BRB
        AntennaGateArea              0.4816 ;
        AntennaPartialMetalArea      2.3500 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2870 LAYER met1 ;
        AntennaDiffArea              0.7350 ;
    END BRB
    PIN GND
    END GND
END RFRDX1
MACRO RF2R1WX2
    PIN WW
        AntennaGateArea              0.2556 ;
        AntennaPartialMetalArea      2.0586 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6398 LAYER met1 ;
    END WW
    PIN WB
        AntennaGateArea              0.1512 ;
        AntennaPartialMetalArea      0.8630 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7380 LAYER met1 ;
    END WB
    PIN R2W
        AntennaGateArea              0.3456 ;
        AntennaPartialMetalArea      1.1014 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0188 LAYER met1 ;
    END R2W
    PIN R2B
        AntennaPartialMetalArea      0.9690 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6066 LAYER met1 ;
        AntennaDiffArea              1.4970 ;
    END R2B
    PIN R1W
        AntennaGateArea              0.3456 ;
        AntennaPartialMetalArea      1.0948 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9864 LAYER met1 ;
    END R1W
    PIN R1B
        AntennaPartialMetalArea      1.0733 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6480 LAYER met1 ;
        AntennaDiffArea              1.4700 ;
    END R1B
    PIN GND
    END GND
END RF2R1WX2
MACRO RF1R1WX2
    PIN WW
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      2.2682 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8522 LAYER met1 ;
    END WW
    PIN WB
        AntennaGateArea              0.1512 ;
        AntennaPartialMetalArea      0.6909 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6228 LAYER met1 ;
    END WB
    PIN RWN
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      1.1068 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9144 LAYER met1 ;
    END RWN
    PIN RW
        AntennaGateArea              0.2160 ;
        AntennaPartialMetalArea      0.7354 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6282 LAYER met1 ;
    END RW
    PIN RB
        AntennaPartialMetalArea      0.6566 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5058 LAYER met1 ;
        AntennaDiffArea              1.3356 ;
    END RB
    PIN GND
    END GND
END RF1R1WX2
MACRO AFCSHCONX4
    PIN S
        AntennaPartialMetalArea      1.5512 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8190 LAYER met1 ;
        AntennaDiffArea              1.4628 ;
    END S
    PIN CS
        AntennaGateArea              0.5832 ;
        AntennaPartialMetalArea      2.4230 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2554 LAYER met1 ;
    END CS
    PIN CO1N
        AntennaPartialMetalArea      2.4898 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6074 LAYER met1 ;
        AntennaDiffArea              3.5424 ;
    END CO1N
    PIN CO0N
        AntennaPartialMetalArea      2.6525 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6992 LAYER met1 ;
        AntennaDiffArea              3.9620 ;
    END CO0N
    PIN CI1
        AntennaGateArea              1.9440 ;
        AntennaPartialMetalArea      2.0362 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4706 LAYER met1 ;
    END CI1
    PIN CI0
        AntennaGateArea              1.8864 ;
        AntennaPartialMetalArea      2.5882 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9710 LAYER met1 ;
    END CI0
    PIN B
        AntennaGateArea              1.5624 ;
        AntennaPartialMetalArea      2.0894 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7334 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              1.0440 ;
        AntennaPartialMetalArea      1.2175 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8640 LAYER met1 ;
    END A
    PIN GND
    END GND
END AFCSHCONX4
MACRO AFCSHCONX2
    PIN S
        AntennaPartialMetalArea      1.3972 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8532 LAYER met1 ;
        AntennaDiffArea              1.3818 ;
    END S
    PIN CS
        AntennaGateArea              0.5832 ;
        AntennaPartialMetalArea      2.4004 LAYER met1 ;
        AntennaPartialMetalSideArea  2.3184 LAYER met1 ;
    END CS
    PIN CO1N
        AntennaPartialMetalArea      1.7256 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1124 LAYER met1 ;
        AntennaDiffArea              2.1394 ;
    END CO1N
    PIN CO0N
        AntennaPartialMetalArea      1.8744 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2870 LAYER met1 ;
        AntennaDiffArea              2.3614 ;
    END CO0N
    PIN CI1
        AntennaGateArea              0.9828 ;
        AntennaPartialMetalArea      1.4682 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0440 LAYER met1 ;
    END CI1
    PIN CI0
        AntennaGateArea              0.9144 ;
        AntennaPartialMetalArea      2.1758 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8036 LAYER met1 ;
    END CI0
    PIN B
        AntennaGateArea              1.4796 ;
        AntennaPartialMetalArea      2.0942 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8054 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              1.0800 ;
        AntennaPartialMetalArea      1.1815 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8280 LAYER met1 ;
    END A
    PIN GND
    END GND
END AFCSHCONX2
MACRO AFCSHCINX4
    PIN S
        AntennaPartialMetalArea      2.1490 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8298 LAYER met1 ;
        AntennaDiffArea              1.3818 ;
    END S
    PIN CS
        AntennaGateArea              0.5832 ;
        AntennaPartialMetalArea      2.3280 LAYER met1 ;
        AntennaPartialMetalSideArea  2.1564 LAYER met1 ;
    END CS
    PIN CO1
        AntennaPartialMetalArea      2.3376 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4940 LAYER met1 ;
        AntennaDiffArea              3.4260 ;
    END CO1
    PIN CO0
        AntennaPartialMetalArea      2.3376 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4940 LAYER met1 ;
        AntennaDiffArea              3.4260 ;
    END CO0
    PIN CI1N
        AntennaGateArea              1.1304 ;
        AntennaPartialMetalArea      1.4652 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0314 LAYER met1 ;
    END CI1N
    PIN CI0N
        AntennaGateArea              1.0728 ;
        AntennaPartialMetalArea      1.7551 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2168 LAYER met1 ;
    END CI0N
    PIN B
        AntennaGateArea              1.5336 ;
        AntennaPartialMetalArea      2.7722 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2590 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      1.2314 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8946 LAYER met1 ;
    END A
    PIN GND
    END GND
END AFCSHCINX4
MACRO AFCSHCINX2
    PIN S
        AntennaPartialMetalArea      2.1490 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8298 LAYER met1 ;
        AntennaDiffArea              1.3818 ;
    END S
    PIN CS
        AntennaGateArea              0.5832 ;
        AntennaPartialMetalArea      2.3280 LAYER met1 ;
        AntennaPartialMetalSideArea  2.1564 LAYER met1 ;
    END CS
    PIN CO1
        AntennaPartialMetalArea      2.3064 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5066 LAYER met1 ;
        AntennaDiffArea              2.5020 ;
    END CO1
    PIN CO0
        AntennaPartialMetalArea      2.2763 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4868 LAYER met1 ;
        AntennaDiffArea              2.4810 ;
    END CO0
    PIN CI1N
        AntennaGateArea              0.6264 ;
        AntennaPartialMetalArea      1.3959 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9252 LAYER met1 ;
    END CI1N
    PIN CI0N
        AntennaGateArea              0.5976 ;
        AntennaPartialMetalArea      1.7383 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1844 LAYER met1 ;
    END CI0N
    PIN B
        AntennaGateArea              1.5336 ;
        AntennaPartialMetalArea      2.7722 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2590 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      1.2314 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8946 LAYER met1 ;
    END A
    PIN GND
    END GND
END AFCSHCINX2
MACRO AHHCONX4
    PIN S
        AntennaPartialMetalArea      1.8907 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2834 LAYER met1 ;
        AntennaDiffArea              1.6440 ;
    END S
    PIN CON
        AntennaPartialMetalArea      2.5654 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2978 LAYER met1 ;
        AntennaDiffArea              3.0538 ;
    END CON
    PIN CI
        AntennaGateArea              1.9764 ;
        AntennaPartialMetalArea      5.1507 LAYER met1 ;
        AntennaPartialMetalSideArea  4.3182 LAYER met1 ;
    END CI
    PIN A
        AntennaGateArea              1.7604 ;
        AntennaPartialMetalArea      2.8128 LAYER met1 ;
        AntennaPartialMetalSideArea  2.0952 LAYER met1 ;
    END A
    PIN GND
    END GND
END AHHCONX4
MACRO AHHCONX2
    PIN S
        AntennaPartialMetalArea      0.9628 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7632 LAYER met1 ;
        AntennaDiffArea              1.6440 ;
    END S
    PIN CON
        AntennaPartialMetalArea      0.9842 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7398 LAYER met1 ;
        AntennaDiffArea              1.3932 ;
    END CON
    PIN CI
        AntennaGateArea              1.3608 ;
        AntennaPartialMetalArea      4.4120 LAYER met1 ;
        AntennaPartialMetalSideArea  3.5082 LAYER met1 ;
    END CI
    PIN A
        AntennaGateArea              1.1448 ;
        AntennaPartialMetalArea      1.8494 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3914 LAYER met1 ;
    END A
    PIN GND
    END GND
END AHHCONX2
MACRO AHHCINX4
    PIN S
    END S
    PIN CO
    END CO
    PIN CIN
    END CIN
    PIN A
    END A
    PIN GND
    END GND
END AHHCINX4
MACRO AHHCINX2
    PIN S
        AntennaPartialMetalArea      0.8612 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6138 LAYER met1 ;
        AntennaDiffArea              1.8912 ;
    END S
    PIN CO
        AntennaPartialMetalArea      0.9200 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6480 LAYER met1 ;
        AntennaDiffArea              1.2960 ;
    END CO
    PIN CIN
        AntennaGateArea              1.4040 ;
        AntennaPartialMetalArea      4.6926 LAYER met1 ;
        AntennaPartialMetalSideArea  3.6972 LAYER met1 ;
    END CIN
    PIN A
        AntennaGateArea              0.7920 ;
        AntennaPartialMetalArea      2.8044 LAYER met1 ;
        AntennaPartialMetalSideArea  2.1978 LAYER met1 ;
    END A
    PIN GND
    END GND
END AHHCINX2
MACRO AFHCONX2
    PIN S
        AntennaPartialMetalArea      2.3218 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8856 LAYER met1 ;
        AntennaDiffArea              1.4308 ;
    END S
    PIN CON
        AntennaPartialMetalArea      2.3558 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4850 LAYER met1 ;
        AntennaDiffArea              2.0358 ;
    END CON
    PIN CI
        AntennaGateArea              1.0584 ;
        AntennaPartialMetalArea      1.3952 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0008 LAYER met1 ;
    END CI
    PIN B
        AntennaGateArea              2.1600 ;
        AntennaPartialMetalArea      2.7358 LAYER met1 ;
        AntennaPartialMetalSideArea  2.1114 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.6886 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5382 LAYER met1 ;
    END A
    PIN GND
    END GND
END AFHCONX2
MACRO AFHCINX2
    PIN S
        AntennaPartialMetalArea      1.8375 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8676 LAYER met1 ;
        AntennaDiffArea              1.3720 ;
    END S
    PIN CO
        AntennaPartialMetalArea      0.9496 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6372 LAYER met1 ;
        AntennaDiffArea              1.5704 ;
    END CO
    PIN CIN
        AntennaGateArea              1.0620 ;
        AntennaPartialMetalArea      1.1322 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8316 LAYER met1 ;
    END CIN
    PIN B
        AntennaGateArea              1.6200 ;
        AntennaPartialMetalArea      3.9508 LAYER met1 ;
        AntennaPartialMetalSideArea  3.7350 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.7022 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6120 LAYER met1 ;
    END A
    PIN GND
    END GND
END AFHCINX2
MACRO CMPR42X2
    PIN S
        AntennaPartialMetalArea      0.8900 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5814 LAYER met1 ;
        AntennaDiffArea              1.4210 ;
    END S
    PIN ICO
        AntennaPartialMetalArea      0.9102 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6246 LAYER met1 ;
        AntennaDiffArea              1.4504 ;
    END ICO
    PIN ICI
        AntennaGateArea              0.4860 ;
        AntennaPartialMetalArea      0.7868 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6228 LAYER met1 ;
    END ICI
    PIN D
        AntennaGateArea              0.9900 ;
        AntennaPartialMetalArea      1.9730 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6326 LAYER met1 ;
    END D
    PIN CO
        AntennaPartialMetalArea      0.7618 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6120 LAYER met1 ;
        AntennaDiffArea              1.1102 ;
    END CO
    PIN C
        AntennaGateArea              0.9036 ;
        AntennaPartialMetalArea      4.8434 LAYER met1 ;
        AntennaPartialMetalSideArea  3.9006 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              1.4688 ;
        AntennaPartialMetalArea      3.8638 LAYER met1 ;
        AntennaPartialMetalSideArea  3.1752 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              1.3140 ;
        AntennaPartialMetalArea      2.9314 LAYER met1 ;
        AntennaPartialMetalSideArea  2.4588 LAYER met1 ;
    END A
    PIN GND
    END GND
END CMPR42X2
MACRO CMPR42X1
    PIN S
        AntennaPartialMetalArea      0.7568 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5004 LAYER met1 ;
        AntennaDiffArea              0.7350 ;
    END S
    PIN ICO
        AntennaPartialMetalArea      0.5784 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4410 LAYER met1 ;
        AntennaDiffArea              0.7350 ;
    END ICO
    PIN ICI
        AntennaGateArea              0.2988 ;
        AntennaPartialMetalArea      0.9824 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8136 LAYER met1 ;
    END ICI
    PIN D
        AntennaGateArea              0.7128 ;
        AntennaPartialMetalArea      1.8930 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7046 LAYER met1 ;
    END D
    PIN CO
        AntennaPartialMetalArea      0.6650 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5094 LAYER met1 ;
        AntennaDiffArea              0.7350 ;
    END CO
    PIN C
        AntennaGateArea              0.5724 ;
        AntennaPartialMetalArea      3.9450 LAYER met1 ;
        AntennaPartialMetalSideArea  3.1428 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.9144 ;
        AntennaPartialMetalArea      3.0272 LAYER met1 ;
        AntennaPartialMetalSideArea  2.7972 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.7884 ;
        AntennaPartialMetalArea      2.3378 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8036 LAYER met1 ;
    END A
    PIN GND
    END GND
END CMPR42X1
MACRO BMXX1
    PIN X2
        AntennaGateArea              0.3384 ;
        AntennaPartialMetalArea      1.0644 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9486 LAYER met1 ;
    END X2
    PIN S
        AntennaGateArea              0.3420 ;
        AntennaPartialMetalArea      0.5493 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4752 LAYER met1 ;
    END S
    PIN PP
        AntennaPartialMetalArea      0.6772 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5148 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END PP
    PIN M1
        AntennaGateArea              0.3132 ;
        AntennaPartialMetalArea      1.6302 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5408 LAYER met1 ;
    END M1
    PIN M0
        AntennaGateArea              0.3132 ;
        AntennaPartialMetalArea      2.0509 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9710 LAYER met1 ;
    END M0
    PIN A
        AntennaGateArea              0.3420 ;
        AntennaPartialMetalArea      0.5292 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4716 LAYER met1 ;
    END A
    PIN GND
    END GND
END BMXX1
MACRO BENCX4
    PIN X2
        AntennaPartialMetalArea      3.1968 LAYER met1 ;
        AntennaPartialMetalSideArea  2.1474 LAYER met1 ;
        AntennaDiffArea              6.4800 ;
    END X2
    PIN S
        AntennaPartialMetalArea      5.2636 LAYER met1 ;
        AntennaPartialMetalSideArea  2.9610 LAYER met1 ;
        AntennaDiffArea              6.4800 ;
    END S
    PIN M2
        AntennaGateArea              0.7740 ;
        AntennaPartialMetalArea      6.9992 LAYER met1 ;
        AntennaPartialMetalSideArea  5.7942 LAYER met1 ;
    END M2
    PIN M1
        AntennaGateArea              2.1996 ;
        AntennaPartialMetalArea      7.1026 LAYER met1 ;
        AntennaPartialMetalSideArea  5.9274 LAYER met1 ;
    END M1
    PIN M0
        AntennaGateArea              2.2032 ;
        AntennaPartialMetalArea      4.8094 LAYER met1 ;
        AntennaPartialMetalSideArea  3.6864 LAYER met1 ;
    END M0
    PIN A
        AntennaPartialMetalArea      6.4201 LAYER met1 ;
        AntennaPartialMetalSideArea  3.2202 LAYER met1 ;
        AntennaDiffArea              6.5040 ;
    END A
    PIN GND
    END GND
END BENCX4
MACRO XOR3X4
    PIN Y
        AntennaPartialMetalArea      1.5125 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7902 LAYER met1 ;
        AntennaDiffArea              1.6200 ;
    END Y
    PIN C
        AntennaGateArea              1.1592 ;
        AntennaPartialMetalArea      2.4296 LAYER met1 ;
        AntennaPartialMetalSideArea  2.3508 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              1.9008 ;
        AntennaPartialMetalArea      4.6734 LAYER met1 ;
        AntennaPartialMetalSideArea  4.3182 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.8267 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5886 LAYER met1 ;
    END A
    PIN GND
    END GND
END XOR3X4
MACRO XOR3X2
    PIN Y
        AntennaPartialMetalArea      0.9712 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6102 LAYER met1 ;
        AntennaDiffArea              1.3945 ;
    END Y
    PIN C
        AntennaGateArea              0.5832 ;
        AntennaPartialMetalArea      1.7282 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6254 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              1.3374 ;
        AntennaPartialMetalArea      3.1526 LAYER met1 ;
        AntennaPartialMetalSideArea  2.9952 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5442 ;
        AntennaPartialMetalArea      0.7716 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5814 LAYER met1 ;
    END A
    PIN GND
    END GND
END XOR3X2
MACRO XNOR3X4
    PIN Y
        AntennaPartialMetalArea      1.5125 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7902 LAYER met1 ;
        AntennaDiffArea              1.6200 ;
    END Y
    PIN C
        AntennaGateArea              1.1664 ;
        AntennaPartialMetalArea      2.4742 LAYER met1 ;
        AntennaPartialMetalSideArea  2.3940 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              1.8972 ;
        AntennaPartialMetalArea      4.6734 LAYER met1 ;
        AntennaPartialMetalSideArea  4.3182 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.8267 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5886 LAYER met1 ;
    END A
    PIN GND
    END GND
END XNOR3X4
MACRO XNOR3X2
    PIN Y
        AntennaPartialMetalArea      0.9672 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6102 LAYER met1 ;
        AntennaDiffArea              1.3945 ;
    END Y
    PIN C
        AntennaGateArea              0.5832 ;
        AntennaPartialMetalArea      1.7876 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6848 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              1.3374 ;
        AntennaPartialMetalArea      3.1526 LAYER met1 ;
        AntennaPartialMetalSideArea  2.9952 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5442 ;
        AntennaPartialMetalArea      0.7281 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5814 LAYER met1 ;
    END A
    PIN GND
    END GND
END XNOR3X2
MACRO AFHCONX4
    PIN S
        AntennaPartialMetalArea      1.7180 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8082 LAYER met1 ;
        AntennaDiffArea              1.4700 ;
    END S
    PIN CON
        AntennaPartialMetalArea      3.3844 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7676 LAYER met1 ;
        AntennaDiffArea              3.0900 ;
    END CON
    PIN CI
        AntennaGateArea              2.1600 ;
        AntennaPartialMetalArea      2.6168 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7316 LAYER met1 ;
    END CI
    PIN B
        AntennaGateArea              2.1600 ;
        AntennaPartialMetalArea      2.7402 LAYER met1 ;
        AntennaPartialMetalSideArea  2.1132 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.6886 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5382 LAYER met1 ;
    END A
    PIN GND
    END GND
END AFHCONX4
MACRO AFHCINX4
    PIN S
        AntennaPartialMetalArea      0.7472 LAYER met1 ;
        AntennaPartialMetalSideArea  0.3852 LAYER met1 ;
        AntennaDiffArea              1.5808 ;
    END S
    PIN CO
        AntennaPartialMetalArea      2.4120 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4004 LAYER met1 ;
        AntennaDiffArea              3.5764 ;
    END CO
    PIN CIN
        AntennaGateArea              2.1600 ;
        AntennaPartialMetalArea      2.6620 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6254 LAYER met1 ;
    END CIN
    PIN B
        AntennaGateArea              1.6200 ;
        AntennaPartialMetalArea      2.1512 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8234 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.8866 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7074 LAYER met1 ;
    END A
    PIN GND
    END GND
END AFHCINX4
MACRO CMPR32X1
    PIN S
        AntennaPartialMetalArea      0.7594 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5598 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END S
    PIN CO
        AntennaPartialMetalArea      0.7574 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5004 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END CO
    PIN C
        AntennaGateArea              0.3816 ;
        AntennaPartialMetalArea      2.0678 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7586 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.6512 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5382 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      1.2278 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8982 LAYER met1 ;
    END A
    PIN GND
    END GND
END CMPR32X1
MACRO CMPR22X1
    PIN S
        AntennaPartialMetalArea      1.0398 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8010 LAYER met1 ;
        AntennaDiffArea              2.3880 ;
    END S
    PIN CO
        AntennaPartialMetalArea      0.7970 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5850 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END CO
    PIN B
        AntennaGateArea              0.8784 ;
        AntennaPartialMetalArea      4.3030 LAYER met1 ;
        AntennaPartialMetalSideArea  3.4434 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.8784 ;
        AntennaPartialMetalArea      1.4427 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0926 LAYER met1 ;
    END A
    PIN GND
    END GND
END CMPR22X1
MACRO BENCX2
    PIN X2
        AntennaPartialMetalArea      1.3881 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0836 LAYER met1 ;
        AntennaDiffArea              3.2400 ;
    END X2
    PIN S
        AntennaPartialMetalArea      2.7016 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3860 LAYER met1 ;
        AntennaDiffArea              3.2400 ;
    END S
    PIN M2
        AntennaGateArea              0.4284 ;
        AntennaPartialMetalArea      4.6511 LAYER met1 ;
        AntennaPartialMetalSideArea  3.8916 LAYER met1 ;
    END M2
    PIN M1
        AntennaGateArea              1.1088 ;
        AntennaPartialMetalArea      4.2592 LAYER met1 ;
        AntennaPartialMetalSideArea  3.6684 LAYER met1 ;
    END M1
    PIN M0
        AntennaGateArea              1.1052 ;
        AntennaPartialMetalArea      3.5899 LAYER met1 ;
        AntennaPartialMetalSideArea  2.8872 LAYER met1 ;
    END M0
    PIN A
        AntennaPartialMetalArea      2.6137 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5588 LAYER met1 ;
        AntennaDiffArea              3.2520 ;
    END A
    PIN GND
    END GND
END BENCX2
MACRO BENCX1
    PIN X2
        AntennaPartialMetalArea      0.7065 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5688 LAYER met1 ;
        AntennaDiffArea              1.6200 ;
    END X2
    PIN S
        AntennaPartialMetalArea      1.1741 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6948 LAYER met1 ;
        AntennaDiffArea              1.6200 ;
    END S
    PIN M2
        AntennaGateArea              0.2844 ;
        AntennaPartialMetalArea      4.3826 LAYER met1 ;
        AntennaPartialMetalSideArea  3.7512 LAYER met1 ;
    END M2
    PIN M1
        AntennaGateArea              0.5580 ;
        AntennaPartialMetalArea      3.9059 LAYER met1 ;
        AntennaPartialMetalSideArea  3.4308 LAYER met1 ;
    END M1
    PIN M0
        AntennaGateArea              0.5544 ;
        AntennaPartialMetalArea      2.8320 LAYER met1 ;
        AntennaPartialMetalSideArea  2.3922 LAYER met1 ;
    END M0
    PIN A
        AntennaPartialMetalArea      1.0454 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7794 LAYER met1 ;
        AntennaDiffArea              1.4998 ;
    END A
    PIN GND
    END GND
END BENCX1
MACRO XOR2XL
    PIN Y
        AntennaPartialMetalArea      1.0516 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6318 LAYER met1 ;
        AntennaDiffArea              0.5582 ;
    END Y
    PIN B
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.8856 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7974 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.3744 ;
        AntennaPartialMetalArea      1.7244 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5570 LAYER met1 ;
    END A
    PIN GND
    END GND
END XOR2XL
MACRO XOR2X4
    PIN Y
        AntennaPartialMetalArea      1.6292 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7344 LAYER met1 ;
        AntennaDiffArea              1.3924 ;
    END Y
    PIN B
        AntennaGateArea              2.3328 ;
        AntennaPartialMetalArea      2.4377 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5642 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              1.2780 ;
        AntennaPartialMetalArea      1.9473 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7280 LAYER met1 ;
    END A
    PIN GND
    END GND
END XOR2X4
MACRO XOR2X2
    PIN Y
        AntennaPartialMetalArea      1.5413 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8208 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Y
    PIN B
        AntennaGateArea              1.1484 ;
        AntennaPartialMetalArea      1.3978 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1862 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.6012 ;
        AntennaPartialMetalArea      1.8650 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5678 LAYER met1 ;
    END A
    PIN GND
    END GND
END XOR2X2
MACRO XOR2X1
    PIN Y
        AntennaPartialMetalArea      1.0516 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6318 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Y
    PIN B
        AntennaGateArea              0.5436 ;
        AntennaPartialMetalArea      0.7084 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6228 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.3456 ;
        AntennaPartialMetalArea      1.7546 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5858 LAYER met1 ;
    END A
    PIN GND
    END GND
END XOR2X1
MACRO XNOR2XL
    PIN Y
        AntennaPartialMetalArea      0.6875 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5058 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END Y
    PIN B
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.5512 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4824 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.3816 ;
        AntennaPartialMetalArea      1.9313 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8396 LAYER met1 ;
    END A
    PIN GND
    END GND
END XNOR2XL
MACRO XNOR2X4
    PIN Y
        AntennaPartialMetalArea      1.6734 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7560 LAYER met1 ;
        AntennaDiffArea              1.3744 ;
    END Y
    PIN B
        AntennaGateArea              2.2032 ;
        AntennaPartialMetalArea      2.1903 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5390 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              1.2420 ;
        AntennaPartialMetalArea      2.0539 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3626 LAYER met1 ;
    END A
    PIN GND
    END GND
END XNOR2X4
MACRO XNOR2X2
    PIN Y
        AntennaPartialMetalArea      1.0826 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6678 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Y
    PIN B
        AntennaGateArea              1.1124 ;
        AntennaPartialMetalArea      1.6281 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2312 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5868 ;
        AntennaPartialMetalArea      2.0944 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7640 LAYER met1 ;
    END A
    PIN GND
    END GND
END XNOR2X2
MACRO XNOR2X1
    PIN Y
        AntennaPartialMetalArea      0.8042 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5688 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Y
    PIN B
        AntennaGateArea              0.4968 ;
        AntennaPartialMetalArea      0.6684 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5364 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.3456 ;
        AntennaPartialMetalArea      2.0722 LAYER met1 ;
        AntennaPartialMetalSideArea  2.0070 LAYER met1 ;
    END A
    PIN GND
    END GND
END XNOR2X1
MACRO TTLATXL
    PIN Q
        AntennaPartialMetalArea      0.6329 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4698 LAYER met1 ;
        AntennaDiffArea              0.4782 ;
    END Q
    PIN OE
        AntennaGateArea              0.1764 ;
        AntennaPartialMetalArea      1.1091 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8676 LAYER met1 ;
    END OE
    PIN G
        AntennaGateArea              0.1260 ;
        AntennaPartialMetalArea      0.6046 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5220 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.6978 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6048 LAYER met1 ;
    END D
    PIN GND
    END GND
END TTLATXL
MACRO TTLATX4
    PIN Q
        AntennaPartialMetalArea      2.7063 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1160 LAYER met1 ;
        AntennaDiffArea              2.8871 ;
    END Q
    PIN OE
        AntennaGateArea              1.1718 ;
        AntennaPartialMetalArea      1.6668 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5120 LAYER met1 ;
    END OE
    PIN G
        AntennaGateArea              0.5292 ;
        AntennaPartialMetalArea      0.7325 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6408 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.9576 ;
        AntennaPartialMetalArea      1.0751 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8856 LAYER met1 ;
    END D
    PIN GND
    END GND
END TTLATX4
MACRO TTLATX2
    PIN Q
        AntennaPartialMetalArea      0.5719 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4284 LAYER met1 ;
        AntennaDiffArea              1.7901 ;
    END Q
    PIN OE
        AntennaGateArea              0.6948 ;
        AntennaPartialMetalArea      1.2752 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0638 LAYER met1 ;
    END OE
    PIN G
        AntennaGateArea              0.3060 ;
        AntennaPartialMetalArea      0.6270 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5436 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.9576 ;
        AntennaPartialMetalArea      1.0893 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9018 LAYER met1 ;
    END D
    PIN GND
    END GND
END TTLATX2
MACRO TTLATX1
    PIN Q
        AntennaPartialMetalArea      1.0143 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7092 LAYER met1 ;
        AntennaDiffArea              1.3357 ;
    END Q
    PIN OE
        AntennaGateArea              0.3420 ;
        AntennaPartialMetalArea      1.1456 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8748 LAYER met1 ;
    END OE
    PIN G
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.6077 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5238 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.5112 ;
        AntennaPartialMetalArea      0.6792 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5796 LAYER met1 ;
    END D
    PIN GND
    END GND
END TTLATX1
MACRO TLATSRXL
    PIN SN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8070 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6444 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.2592 ;
        AntennaPartialMetalArea      1.2954 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2024 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.6836 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4914 LAYER met1 ;
        AntennaDiffArea              0.5853 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6496 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4932 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END Q
    PIN G
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7640 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6786 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.7373 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6588 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATSRXL
MACRO TLATSRX4
    PIN SN
        AntennaGateArea              0.5292 ;
        AntennaPartialMetalArea      0.6580 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5526 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.8640 ;
        AntennaPartialMetalArea      1.9980 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9188 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.1098 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5562 LAYER met1 ;
        AntennaDiffArea              1.4292 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8924 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4734 LAYER met1 ;
        AntennaDiffArea              1.4292 ;
    END Q
    PIN G
        AntennaGateArea              0.3060 ;
        AntennaPartialMetalArea      0.6578 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5850 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.8424 ;
        AntennaPartialMetalArea      2.0456 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9134 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATSRX4
MACRO TLATSRX2
    PIN SN
        AntennaGateArea              0.2988 ;
        AntennaPartialMetalArea      0.6558 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5544 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.4716 ;
        AntennaPartialMetalArea      1.2702 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1736 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.6629 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4590 LAYER met1 ;
        AntennaDiffArea              1.2077 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8300 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6462 LAYER met1 ;
        AntennaDiffArea              1.1699 ;
    END Q
    PIN G
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.7718 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6984 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.4212 ;
        AntennaPartialMetalArea      0.6504 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5814 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATSRX2
MACRO TLATSRX1
    PIN SN
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.7472 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6156 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.3060 ;
        AntennaPartialMetalArea      1.2567 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2150 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.6644 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4824 LAYER met1 ;
        AntennaDiffArea              0.7740 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.5919 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4824 LAYER met1 ;
        AntennaDiffArea              0.8044 ;
    END Q
    PIN G
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.7325 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6534 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.6892 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6390 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATSRX1
MACRO TLATSXL
    PIN SN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7332 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6408 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      0.6023 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4752 LAYER met1 ;
        AntennaDiffArea              0.5674 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.5847 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4770 LAYER met1 ;
        AntennaDiffArea              0.5950 ;
    END Q
    PIN G
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7994 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7452 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.1836 ;
        AntennaPartialMetalArea      0.7165 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6498 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATSXL
MACRO TLATSX4
    PIN SN
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.6509 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5922 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      1.1027 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5544 LAYER met1 ;
        AntennaDiffArea              1.4382 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8924 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4734 LAYER met1 ;
        AntennaDiffArea              1.4382 ;
    END Q
    PIN G
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.8140 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7452 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.7344 ;
        AntennaPartialMetalArea      1.4566 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2906 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATSX4
MACRO TLATSX2
    PIN SN
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.6567 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6012 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      0.8806 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6768 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6636 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5166 LAYER met1 ;
        AntennaDiffArea              1.0823 ;
    END Q
    PIN G
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.8126 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7668 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.4104 ;
        AntennaPartialMetalArea      0.7273 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6444 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATSX2
MACRO TLATSX1
    PIN SN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6853 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5976 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      0.6608 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4806 LAYER met1 ;
        AntennaDiffArea              0.7740 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.5903 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4644 LAYER met1 ;
        AntennaDiffArea              0.8044 ;
    END Q
    PIN G
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.8976 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7416 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.2304 ;
        AntennaPartialMetalArea      0.7056 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6246 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATSX1
MACRO TLATRXL
    PIN RN
        AntennaGateArea              0.2340 ;
        AntennaPartialMetalArea      1.7836 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5606 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.6806 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5076 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.2033 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9450 LAYER met1 ;
        AntennaDiffArea              0.5896 ;
    END Q
    PIN G
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6404 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5616 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.9709 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9054 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATRXL
MACRO TLATRX4
    PIN RN
        AntennaGateArea              0.5040 ;
        AntennaPartialMetalArea      1.6613 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5660 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.8520 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4374 LAYER met1 ;
        AntennaDiffArea              1.7232 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.0824 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4788 LAYER met1 ;
        AntennaDiffArea              1.6200 ;
    END Q
    PIN G
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.7866 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6804 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.7992 ;
        AntennaPartialMetalArea      1.3750 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1448 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATRX4
MACRO TLATRX2
    PIN RN
        AntennaGateArea              0.3420 ;
        AntennaPartialMetalArea      1.7966 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6020 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.8854 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6336 LAYER met1 ;
        AntennaDiffArea              1.2728 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.7327 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5904 LAYER met1 ;
        AntennaDiffArea              1.1018 ;
    END Q
    PIN G
        AntennaGateArea              0.1692 ;
        AntennaPartialMetalArea      0.6455 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5598 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.4212 ;
        AntennaPartialMetalArea      0.7581 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6858 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATRX2
MACRO TLATRX1
    PIN RN
        AntennaGateArea              0.2556 ;
        AntennaPartialMetalArea      1.8556 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6722 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.6971 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4896 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.2465 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9774 LAYER met1 ;
        AntennaDiffArea              0.7680 ;
    END Q
    PIN G
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.6528 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5616 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      1.1123 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8856 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATRX1
MACRO TLATNSRXL
    PIN SN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7898 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7020 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.2592 ;
        AntennaPartialMetalArea      1.2394 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1988 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.6848 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4914 LAYER met1 ;
        AntennaDiffArea              0.5853 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6039 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4914 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END Q
    PIN GN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9305 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8514 LAYER met1 ;
    END GN
    PIN D
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.7666 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6606 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATNSRXL
MACRO TLATNSRX4
    PIN SN
        AntennaGateArea              0.5292 ;
        AntennaPartialMetalArea      0.6356 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5364 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.8640 ;
        AntennaPartialMetalArea      1.9660 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9008 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.1205 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5544 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8924 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4734 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END Q
    PIN GN
        AntennaGateArea              0.3060 ;
        AntennaPartialMetalArea      0.6640 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5940 LAYER met1 ;
    END GN
    PIN D
        AntennaGateArea              0.8424 ;
        AntennaPartialMetalArea      2.0505 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9170 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATNSRX4
MACRO TLATNSRX2
    PIN SN
        AntennaGateArea              0.2988 ;
        AntennaPartialMetalArea      0.8604 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7650 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.4716 ;
        AntennaPartialMetalArea      1.1946 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1160 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.6323 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4482 LAYER met1 ;
        AntennaDiffArea              1.2758 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.7576 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5868 LAYER met1 ;
        AntennaDiffArea              1.2438 ;
    END Q
    PIN GN
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.7713 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6966 LAYER met1 ;
    END GN
    PIN D
        AntennaGateArea              0.4212 ;
        AntennaPartialMetalArea      0.6043 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5148 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATNSRX2
MACRO TLATNSRX1
    PIN SN
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.9532 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7254 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.3060 ;
        AntennaPartialMetalArea      1.2339 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1952 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.6606 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4824 LAYER met1 ;
        AntennaDiffArea              0.7740 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.5919 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4824 LAYER met1 ;
        AntennaDiffArea              0.7986 ;
    END Q
    PIN GN
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.8132 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7326 LAYER met1 ;
    END GN
    PIN D
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.6862 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6390 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATNSRX1
MACRO TLATNSXL
    PIN SN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7134 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6120 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      0.6023 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4752 LAYER met1 ;
        AntennaDiffArea              0.5674 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.5847 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4770 LAYER met1 ;
        AntennaDiffArea              0.6046 ;
    END Q
    PIN GN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8461 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7956 LAYER met1 ;
    END GN
    PIN D
        AntennaGateArea              0.1836 ;
        AntennaPartialMetalArea      0.7372 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6516 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATNSXL
MACRO TLATNSX4
    PIN SN
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.6345 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5598 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      0.9843 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5544 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8966 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4734 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END Q
    PIN GN
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.9092 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8370 LAYER met1 ;
    END GN
    PIN D
        AntennaGateArea              0.7344 ;
        AntennaPartialMetalArea      1.4519 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2780 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATNSX4
MACRO TLATNSX2
    PIN SN
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.6686 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5832 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      0.8690 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6930 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.7218 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5616 LAYER met1 ;
        AntennaDiffArea              1.1844 ;
    END Q
    PIN GN
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.6368 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5886 LAYER met1 ;
    END GN
    PIN D
        AntennaGateArea              0.4104 ;
        AntennaPartialMetalArea      0.6104 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5400 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATNSX2
MACRO TLATNSX1
    PIN SN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6748 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5832 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      0.6568 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4806 LAYER met1 ;
        AntennaDiffArea              0.7350 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.5812 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4752 LAYER met1 ;
        AntennaDiffArea              0.7542 ;
    END Q
    PIN GN
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.7437 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6966 LAYER met1 ;
    END GN
    PIN D
        AntennaGateArea              0.2304 ;
        AntennaPartialMetalArea      0.7445 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6714 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATNSX1
MACRO TLATNRXL
    PIN RN
        AntennaGateArea              0.2376 ;
        AntennaPartialMetalArea      1.7666 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5876 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.7204 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5220 LAYER met1 ;
        AntennaDiffArea              0.5484 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.2447 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9612 LAYER met1 ;
        AntennaDiffArea              0.5484 ;
    END Q
    PIN GN
        AntennaGateArea              0.1332 ;
        AntennaPartialMetalArea      0.6708 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5274 LAYER met1 ;
    END GN
    PIN D
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.7756 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7056 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATNRXL
MACRO TLATNRX4
    PIN RN
        AntennaGateArea              0.4824 ;
        AntennaPartialMetalArea      1.6532 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5840 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.8338 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4482 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.0428 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5760 LAYER met1 ;
        AntennaDiffArea              1.7400 ;
    END Q
    PIN GN
        AntennaGateArea              0.2628 ;
        AntennaPartialMetalArea      0.7544 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6624 LAYER met1 ;
    END GN
    PIN D
        AntennaGateArea              0.7776 ;
        AntennaPartialMetalArea      1.4264 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1826 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATNRX4
MACRO TLATNRX2
    PIN RN
        AntennaGateArea              0.3420 ;
        AntennaPartialMetalArea      1.8664 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6074 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.0934 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6822 LAYER met1 ;
        AntennaDiffArea              1.6320 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8855 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6678 LAYER met1 ;
        AntennaDiffArea              1.1652 ;
    END Q
    PIN GN
        AntennaGateArea              0.1620 ;
        AntennaPartialMetalArea      0.7220 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5814 LAYER met1 ;
    END GN
    PIN D
        AntennaGateArea              0.4212 ;
        AntennaPartialMetalArea      0.8129 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7236 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATNRX2
MACRO TLATNRX1
    PIN RN
        AntennaGateArea              0.2556 ;
        AntennaPartialMetalArea      1.7696 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5912 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.6568 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4896 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.2447 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9612 LAYER met1 ;
        AntennaDiffArea              0.8040 ;
    END Q
    PIN GN
        AntennaGateArea              0.1332 ;
        AntennaPartialMetalArea      0.6708 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5274 LAYER met1 ;
    END GN
    PIN D
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      0.7261 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6624 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATNRX1
MACRO TLATNXL
    PIN QN
        AntennaPartialMetalArea      0.6958 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5184 LAYER met1 ;
        AntennaDiffArea              0.5938 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.3244 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0080 LAYER met1 ;
        AntennaDiffArea              0.6130 ;
    END Q
    PIN GN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6698 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5472 LAYER met1 ;
    END GN
    PIN D
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7670 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6714 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATNXL
MACRO TLATNX4
    PIN QN
        AntennaPartialMetalArea      0.8854 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4518 LAYER met1 ;
        AntennaDiffArea              1.4574 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8800 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4806 LAYER met1 ;
        AntennaDiffArea              1.4232 ;
    END Q
    PIN GN
        AntennaGateArea              0.3420 ;
        AntennaPartialMetalArea      0.7368 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5850 LAYER met1 ;
    END GN
    PIN D
        AntennaGateArea              1.0800 ;
        AntennaPartialMetalArea      2.4818 LAYER met1 ;
        AntennaPartialMetalSideArea  2.0124 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATNX4
MACRO TLATNX2
    PIN QN
        AntennaPartialMetalArea      1.1017 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6606 LAYER met1 ;
        AntennaDiffArea              1.6560 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.9569 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6930 LAYER met1 ;
        AntennaDiffArea              1.2158 ;
    END Q
    PIN GN
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.7042 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5688 LAYER met1 ;
    END GN
    PIN D
        AntennaGateArea              0.5184 ;
        AntennaPartialMetalArea      0.7002 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6048 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATNX2
MACRO TLATNX1
    PIN QN
        AntennaPartialMetalArea      0.6876 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4896 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.3300 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0062 LAYER met1 ;
        AntennaDiffArea              0.8040 ;
    END Q
    PIN GN
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.6738 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5562 LAYER met1 ;
    END GN
    PIN D
        AntennaGateArea              0.3024 ;
        AntennaPartialMetalArea      0.7360 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6678 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATNX1
MACRO TLATXL
    PIN QN
        AntennaPartialMetalArea      0.6900 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5220 LAYER met1 ;
        AntennaDiffArea              0.5938 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.2437 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9558 LAYER met1 ;
        AntennaDiffArea              0.6322 ;
    END Q
    PIN G
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7272 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5760 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.8928 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7650 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATXL
MACRO TLATX4
    PIN QN
        AntennaPartialMetalArea      0.8854 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4518 LAYER met1 ;
        AntennaDiffArea              1.4574 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8800 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4806 LAYER met1 ;
        AntennaDiffArea              1.4232 ;
    END Q
    PIN G
        AntennaGateArea              0.3420 ;
        AntennaPartialMetalArea      0.7653 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5904 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              1.0800 ;
        AntennaPartialMetalArea      2.4818 LAYER met1 ;
        AntennaPartialMetalSideArea  2.0124 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATX4
MACRO TLATX2
    PIN QN
        AntennaPartialMetalArea      1.3260 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7344 LAYER met1 ;
        AntennaDiffArea              1.6800 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.7824 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6012 LAYER met1 ;
        AntennaDiffArea              1.1948 ;
    END Q
    PIN G
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.7206 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5868 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.5184 ;
        AntennaPartialMetalArea      0.6871 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5922 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATX2
MACRO TLATX1
    PIN QN
        AntennaPartialMetalArea      0.6568 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4896 LAYER met1 ;
        AntennaDiffArea              0.8400 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.3327 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0224 LAYER met1 ;
        AntennaDiffArea              0.8040 ;
    END Q
    PIN G
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.6919 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5634 LAYER met1 ;
    END G
    PIN D
        AntennaGateArea              0.3132 ;
        AntennaPartialMetalArea      0.7370 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6696 LAYER met1 ;
    END D
    PIN GND
    END GND
END TLATX1
MACRO TIELO
    PIN Y
        AntennaPartialMetalArea      0.2760 LAYER met1 ;
        AntennaPartialMetalSideArea  0.1908 LAYER met1 ;
        AntennaDiffArea              0.5712 ;
    END Y
    PIN GND
    END GND
END TIELO
MACRO TIEHI
    PIN Y
        AntennaPartialMetalArea      0.2661 LAYER met1 ;
        AntennaPartialMetalSideArea  0.2160 LAYER met1 ;
        AntennaDiffArea              0.4739 ;
    END Y
    PIN GND
    END GND
END TIEHI
MACRO TBUFIXL
    PIN Y
        AntennaPartialMetalArea      1.2486 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7344 LAYER met1 ;
        AntennaDiffArea              1.1172 ;
    END Y
    PIN OE
        AntennaGateArea              0.2808 ;
        AntennaPartialMetalArea      1.2227 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1340 LAYER met1 ;
    END OE
    PIN A
        AntennaGateArea              0.3780 ;
        AntennaPartialMetalArea      0.6498 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5904 LAYER met1 ;
    END A
    PIN GND
    END GND
END TBUFIXL
MACRO TBUFIX8
    PIN Y
        AntennaPartialMetalArea      4.4514 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1250 LAYER met1 ;
        AntennaDiffArea              3.4730 ;
    END Y
    PIN OE
        AntennaGateArea              0.4788 ;
        AntennaPartialMetalArea      1.6056 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4328 LAYER met1 ;
    END OE
    PIN A
        AntennaGateArea              0.3420 ;
        AntennaPartialMetalArea      0.6633 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6030 LAYER met1 ;
    END A
    PIN GND
    END GND
END TBUFIX8
MACRO TBUFIX4
    PIN Y
        AntennaPartialMetalArea      1.2832 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5868 LAYER met1 ;
        AntennaDiffArea              1.6374 ;
    END Y
    PIN OE
        AntennaGateArea              0.2952 ;
        AntennaPartialMetalArea      1.6274 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4742 LAYER met1 ;
    END OE
    PIN A
        AntennaGateArea              0.1692 ;
        AntennaPartialMetalArea      1.3846 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1790 LAYER met1 ;
    END A
    PIN GND
    END GND
END TBUFIX4
MACRO TBUFIX3
    PIN Y
        AntennaPartialMetalArea      1.2639 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7182 LAYER met1 ;
        AntennaDiffArea              1.3108 ;
    END Y
    PIN OE
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      1.6196 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5084 LAYER met1 ;
    END OE
    PIN A
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      1.3514 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1844 LAYER met1 ;
    END A
    PIN GND
    END GND
END TBUFIX3
MACRO TBUFIX2
    PIN Y
        AntennaPartialMetalArea      1.4486 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0224 LAYER met1 ;
        AntennaDiffArea              1.1400 ;
    END Y
    PIN OE
        AntennaGateArea              0.4572 ;
        AntennaPartialMetalArea      1.8196 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5138 LAYER met1 ;
    END OE
    PIN A
        AntennaGateArea              0.7200 ;
        AntennaPartialMetalArea      1.7148 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4706 LAYER met1 ;
    END A
    PIN GND
    END GND
END TBUFIX2
MACRO TBUFIX20
    PIN Y
        AntennaPartialMetalArea      12.0036 LAYER met1 ;
        AntennaPartialMetalSideArea  2.6154 LAYER met1 ;
        AntennaDiffArea              8.5962 ;
    END Y
    PIN OE
        AntennaGateArea              1.1616 ;
        AntennaPartialMetalArea      1.7742 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6560 LAYER met1 ;
    END OE
    PIN A
        AntennaGateArea              0.8460 ;
        AntennaPartialMetalArea      1.2353 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8946 LAYER met1 ;
    END A
    PIN GND
    END GND
END TBUFIX20
MACRO TBUFIX1
    PIN Y
        AntennaPartialMetalArea      1.2706 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7866 LAYER met1 ;
        AntennaDiffArea              1.1560 ;
    END Y
    PIN OE
        AntennaGateArea              0.2736 ;
        AntennaPartialMetalArea      1.2079 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0386 LAYER met1 ;
    END OE
    PIN A
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7768 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6768 LAYER met1 ;
    END A
    PIN GND
    END GND
END TBUFIX1
MACRO TBUFIX16
    PIN Y
        AntennaPartialMetalArea      9.9108 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2032 LAYER met1 ;
        AntennaDiffArea              6.8588 ;
    END Y
    PIN OE
        AntennaGateArea              0.9540 ;
        AntennaPartialMetalArea      1.8038 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7136 LAYER met1 ;
    END OE
    PIN A
        AntennaGateArea              0.6732 ;
        AntennaPartialMetalArea      1.2772 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9468 LAYER met1 ;
    END A
    PIN GND
    END GND
END TBUFIX16
MACRO TBUFIX12
    PIN Y
        AntennaPartialMetalArea      6.7022 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5570 LAYER met1 ;
        AntennaDiffArea              5.2020 ;
    END Y
    PIN OE
        AntennaGateArea              0.7282 ;
        AntennaPartialMetalArea      1.7976 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6740 LAYER met1 ;
    END OE
    PIN A
        AntennaGateArea              0.5148 ;
        AntennaPartialMetalArea      0.6435 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5832 LAYER met1 ;
    END A
    PIN GND
    END GND
END TBUFIX12
MACRO TBUFXL
    PIN Y
        AntennaPartialMetalArea      1.2840 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6498 LAYER met1 ;
        AntennaDiffArea              0.5906 ;
    END Y
    PIN OE
        AntennaGateArea              0.2376 ;
        AntennaPartialMetalArea      1.2437 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1520 LAYER met1 ;
    END OE
    PIN A
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8940 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8100 LAYER met1 ;
    END A
    PIN GND
    END GND
END TBUFXL
MACRO TBUFX8
    PIN Y
        AntennaPartialMetalArea      5.5809 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1340 LAYER met1 ;
        AntennaDiffArea              3.2619 ;
    END Y
    PIN OE
        AntennaGateArea              0.4788 ;
        AntennaPartialMetalArea      1.2106 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1178 LAYER met1 ;
    END OE
    PIN A
        AntennaGateArea              0.8496 ;
        AntennaPartialMetalArea      1.9687 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6398 LAYER met1 ;
    END A
    PIN GND
    END GND
END TBUFX8
MACRO TBUFX4
    PIN Y
        AntennaPartialMetalArea      1.4768 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7560 LAYER met1 ;
        AntennaDiffArea              1.7400 ;
    END Y
    PIN OE
        AntennaGateArea              0.3024 ;
        AntennaPartialMetalArea      1.7217 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6416 LAYER met1 ;
    END OE
    PIN A
        AntennaGateArea              0.4320 ;
        AntennaPartialMetalArea      0.8504 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7524 LAYER met1 ;
    END A
    PIN GND
    END GND
END TBUFX4
MACRO TBUFX3
    PIN Y
        AntennaPartialMetalArea      1.6500 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7146 LAYER met1 ;
        AntennaDiffArea              1.1596 ;
    END Y
    PIN OE
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      1.2467 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1718 LAYER met1 ;
    END OE
    PIN A
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      0.7706 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7236 LAYER met1 ;
    END A
    PIN GND
    END GND
END TBUFX3
MACRO TBUFX2
    PIN Y
        AntennaPartialMetalArea      0.8108 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5904 LAYER met1 ;
        AntennaDiffArea              1.2267 ;
    END Y
    PIN OE
        AntennaGateArea              0.2592 ;
        AntennaPartialMetalArea      1.3038 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1916 LAYER met1 ;
    END OE
    PIN A
        AntennaGateArea              0.2160 ;
        AntennaPartialMetalArea      0.8886 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7938 LAYER met1 ;
    END A
    PIN GND
    END GND
END TBUFX2
MACRO TBUFX20
    PIN Y
        AntennaPartialMetalArea      11.6440 LAYER met1 ;
        AntennaPartialMetalSideArea  2.4318 LAYER met1 ;
        AntennaDiffArea              7.5274 ;
    END Y
    PIN OE
        AntennaGateArea              1.1916 ;
        AntennaPartialMetalArea      2.1530 LAYER met1 ;
        AntennaPartialMetalSideArea  2.0340 LAYER met1 ;
    END OE
    PIN A
        AntennaGateArea              2.2400 ;
        AntennaPartialMetalArea      2.7381 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8252 LAYER met1 ;
    END A
    PIN GND
    END GND
END TBUFX20
MACRO TBUFX1
    PIN Y
        AntennaPartialMetalArea      1.2518 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6174 LAYER met1 ;
        AntennaDiffArea              0.8220 ;
    END Y
    PIN OE
        AntennaGateArea              0.2592 ;
        AntennaPartialMetalArea      1.2537 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1880 LAYER met1 ;
    END OE
    PIN A
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9468 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8478 LAYER met1 ;
    END A
    PIN GND
    END GND
END TBUFX1
MACRO TBUFX16
    PIN Y
        AntennaPartialMetalArea      10.0382 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9278 LAYER met1 ;
        AntennaDiffArea              5.8782 ;
    END Y
    PIN OE
        AntennaGateArea              0.9576 ;
        AntennaPartialMetalArea      1.6218 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5084 LAYER met1 ;
    END OE
    PIN A
        AntennaGateArea              1.7604 ;
        AntennaPartialMetalArea      1.7422 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2582 LAYER met1 ;
    END A
    PIN GND
    END GND
END TBUFX16
MACRO TBUFX12
    PIN Y
        AntennaPartialMetalArea      6.9073 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5606 LAYER met1 ;
        AntennaDiffArea              5.0592 ;
    END Y
    PIN OE
        AntennaGateArea              0.7200 ;
        AntennaPartialMetalArea      1.6366 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3770 LAYER met1 ;
    END OE
    PIN A
        AntennaGateArea              1.3524 ;
        AntennaPartialMetalArea      1.8279 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3284 LAYER met1 ;
    END A
    PIN GND
    END GND
END TBUFX12
MACRO SEDFFTRXL
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7830 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6930 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2844 ;
        AntennaPartialMetalArea      0.9380 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8226 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      1.0502 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9774 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.2134 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9108 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.7569 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5400 LAYER met1 ;
        AntennaDiffArea              0.6600 ;
    END Q
    PIN E
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.5360 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4734 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.5846 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5040 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.5688 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4932 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SEDFFTRXL
MACRO SEDFFTRX4
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7326 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6426 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2844 ;
        AntennaPartialMetalArea      0.9168 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7668 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      1.0358 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9630 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.9520 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4824 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.3414 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7956 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END Q
    PIN E
        AntennaGateArea              0.1332 ;
        AntennaPartialMetalArea      0.5360 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4734 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.2160 ;
        AntennaPartialMetalArea      0.5646 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4950 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.5381 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4752 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SEDFFTRX4
MACRO SEDFFTRX2
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7686 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6588 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2844 ;
        AntennaPartialMetalArea      0.9086 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7650 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      1.0358 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9630 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.5778 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4554 LAYER met1 ;
        AntennaDiffArea              1.2401 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8040 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5886 LAYER met1 ;
        AntennaDiffArea              1.2227 ;
    END Q
    PIN E
        AntennaGateArea              0.1332 ;
        AntennaPartialMetalArea      0.5716 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4896 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.2160 ;
        AntennaPartialMetalArea      0.5660 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4950 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.5629 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4896 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SEDFFTRX2
MACRO SEDFFTRX1
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7294 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6426 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2844 ;
        AntennaPartialMetalArea      0.9112 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7668 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.9999 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9252 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.7352 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5472 LAYER met1 ;
        AntennaDiffArea              0.7372 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.7622 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5616 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN E
        AntennaGateArea              0.1332 ;
        AntennaPartialMetalArea      0.5636 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4860 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.2160 ;
        AntennaPartialMetalArea      0.5660 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4950 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.5399 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4770 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SEDFFTRX1
MACRO SEDFFHQXL
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8131 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7164 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6857 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5598 LAYER met1 ;
    END SE
    PIN Q
        AntennaPartialMetalArea      0.8505 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6282 LAYER met1 ;
        AntennaDiffArea              0.5200 ;
    END Q
    PIN E
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7088 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6426 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.5947 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5310 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6904 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5724 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SEDFFHQXL
MACRO SEDFFHQX4
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8633 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7218 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6931 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5688 LAYER met1 ;
    END SE
    PIN Q
        AntennaPartialMetalArea      1.7604 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8226 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END Q
    PIN E
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6958 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6282 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.6534 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5580 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.5220 ;
        AntennaPartialMetalArea      0.7388 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5904 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SEDFFHQX4
MACRO SEDFFHQX2
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8368 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7200 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6931 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5688 LAYER met1 ;
    END SE
    PIN Q
        AntennaPartialMetalArea      0.8420 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5616 LAYER met1 ;
        AntennaDiffArea              1.2455 ;
    END Q
    PIN E
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7037 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6282 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.6516 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5580 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.3420 ;
        AntennaPartialMetalArea      0.7430 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6012 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SEDFFHQX2
MACRO SEDFFHQX1
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8596 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7218 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6965 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5706 LAYER met1 ;
    END SE
    PIN Q
        AntennaPartialMetalArea      0.8220 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5958 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN E
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7035 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6534 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.6602 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5850 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.6553 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5454 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SEDFFHQX1
MACRO SEDFFXL
    PIN SI
        AntennaGateArea              0.1260 ;
        AntennaPartialMetalArea      0.7612 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6912 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      1.6028 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4940 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      0.6277 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4392 LAYER met1 ;
        AntennaDiffArea              0.6422 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.2110 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9054 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END Q
    PIN E
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      2.6602 LAYER met1 ;
        AntennaPartialMetalSideArea  2.5524 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.1260 ;
        AntennaPartialMetalArea      0.8428 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7776 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1260 ;
        AntennaPartialMetalArea      0.7143 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6336 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SEDFFXL
MACRO SEDFFX4
    PIN SI
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.7286 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6606 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.3960 ;
        AntennaPartialMetalArea      1.9520 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8432 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      0.8644 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4428 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.9444 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4788 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END Q
    PIN E
        AntennaGateArea              0.3744 ;
        AntennaPartialMetalArea      2.6656 LAYER met1 ;
        AntennaPartialMetalSideArea  2.5578 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.2376 ;
        AntennaPartialMetalArea      0.7839 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7236 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.5220 ;
        AntennaPartialMetalArea      0.8686 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7290 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SEDFFX4
MACRO SEDFFX2
    PIN SI
        AntennaGateArea              0.1404 ;
        AntennaPartialMetalArea      0.7592 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6876 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2844 ;
        AntennaPartialMetalArea      1.8890 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8306 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      0.9222 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6048 LAYER met1 ;
        AntennaDiffArea              1.4350 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6727 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4680 LAYER met1 ;
        AntennaDiffArea              1.1894 ;
    END Q
    PIN E
        AntennaGateArea              0.2664 ;
        AntennaPartialMetalArea      2.6593 LAYER met1 ;
        AntennaPartialMetalSideArea  2.5524 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.1404 ;
        AntennaPartialMetalArea      0.8268 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7812 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.3060 ;
        AntennaPartialMetalArea      0.5545 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4932 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SEDFFX2
MACRO SEDFFX1
    PIN SI
        AntennaGateArea              0.1008 ;
        AntennaPartialMetalArea      0.8116 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7416 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2340 ;
        AntennaPartialMetalArea      1.8332 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7280 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      0.6874 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5004 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.2710 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9540 LAYER met1 ;
        AntennaDiffArea              0.7530 ;
    END Q
    PIN E
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      2.6845 LAYER met1 ;
        AntennaPartialMetalSideArea  2.5776 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.1008 ;
        AntennaPartialMetalArea      0.8824 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8082 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2052 ;
        AntennaPartialMetalArea      0.6816 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6192 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SEDFFX1
MACRO SDFFTRXL
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9629 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9090 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.3024 ;
        AntennaPartialMetalArea      1.8499 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5894 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.1944 ;
        AntennaPartialMetalArea      0.9604 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8694 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.9007 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5904 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.4019 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0188 LAYER met1 ;
        AntennaDiffArea              0.5628 ;
    END Q
    PIN D
        AntennaGateArea              0.1944 ;
        AntennaPartialMetalArea      1.1128 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0692 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6606 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5598 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFTRXL
MACRO SDFFTRX4
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9573 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8694 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      2.3861 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9134 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.2412 ;
        AntennaPartialMetalArea      1.5586 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2996 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.1107 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4824 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.0259 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4554 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END Q
    PIN D
        AntennaGateArea              0.2412 ;
        AntennaPartialMetalArea      0.8285 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7380 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.5040 ;
        AntennaPartialMetalArea      0.5893 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4968 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFTRX4
MACRO SDFFTRX2
    PIN SI
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.8883 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7614 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2664 ;
        AntennaPartialMetalArea      1.6967 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6074 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.8420 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7830 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.0452 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6966 LAYER met1 ;
        AntennaDiffArea              1.5780 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.7842 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5652 LAYER met1 ;
        AntennaDiffArea              1.2292 ;
    END Q
    PIN D
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      1.0271 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9540 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      0.6914 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6102 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFTRX2
MACRO SDFFTRX1
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9400 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8874 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2376 ;
        AntennaPartialMetalArea      1.7963 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5786 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      1.0644 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9378 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.8390 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5688 LAYER met1 ;
        AntennaDiffArea              0.7860 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.4744 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0602 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN D
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      1.0938 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0350 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2016 ;
        AntennaPartialMetalArea      0.6910 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5580 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFTRX1
MACRO SDFFSRHQXL
    PIN SN
        AntennaGateArea              0.4968 ;
        AntennaPartialMetalArea      5.7438 LAYER met1 ;
        AntennaPartialMetalSideArea  4.5360 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6500 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5814 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.3024 ;
        AntennaPartialMetalArea      2.4678 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2446 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7248 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6660 LAYER met1 ;
    END RN
    PIN Q
        AntennaPartialMetalArea      1.1820 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8586 LAYER met1 ;
        AntennaDiffArea              0.7760 ;
    END Q
    PIN D
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.9849 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8568 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8475 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7686 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFSRHQXL
MACRO SDFFSRHQX4
    PIN SN
        AntennaGateArea              1.7562 ;
        AntennaPartialMetalArea      7.6488 LAYER met1 ;
        AntennaPartialMetalSideArea  5.6790 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6912 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6030 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.3672 ;
        AntennaPartialMetalArea      2.5492 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2968 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.8136 ;
        AntennaPartialMetalArea      1.3250 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9828 LAYER met1 ;
    END RN
    PIN Q
        AntennaPartialMetalArea      3.6404 LAYER met1 ;
        AntennaPartialMetalSideArea  2.3238 LAYER met1 ;
        AntennaDiffArea              4.8883 ;
    END Q
    PIN D
        AntennaGateArea              0.3096 ;
        AntennaPartialMetalArea      0.8120 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6930 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.5148 ;
        AntennaPartialMetalArea      0.7424 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5850 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFSRHQX4
MACRO SDFFSRHQX2
    PIN SN
        AntennaGateArea              0.9720 ;
        AntennaPartialMetalArea      6.5031 LAYER met1 ;
        AntennaPartialMetalSideArea  5.0508 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6486 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5814 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2916 ;
        AntennaPartialMetalArea      2.4776 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2572 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.4428 ;
        AntennaPartialMetalArea      0.6858 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5796 LAYER met1 ;
    END RN
    PIN Q
        AntennaPartialMetalArea      1.8539 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2888 LAYER met1 ;
        AntennaDiffArea              2.5965 ;
    END Q
    PIN D
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.7647 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5976 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.3060 ;
        AntennaPartialMetalArea      0.6107 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5238 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFSRHQX2
MACRO SDFFSRHQX1
    PIN SN
        AntennaGateArea              0.5688 ;
        AntennaPartialMetalArea      5.7114 LAYER met1 ;
        AntennaPartialMetalSideArea  4.5036 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6500 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5814 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      2.5020 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2788 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7116 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6462 LAYER met1 ;
    END RN
    PIN Q
        AntennaPartialMetalArea      1.1464 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8802 LAYER met1 ;
        AntennaDiffArea              1.1060 ;
    END Q
    PIN D
        AntennaGateArea              0.1224 ;
        AntennaPartialMetalArea      0.6409 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5796 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2052 ;
        AntennaPartialMetalArea      0.5921 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5058 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFSRHQX1
MACRO SDFFSRXL
    PIN SN
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      3.2649 LAYER met1 ;
        AntennaPartialMetalSideArea  2.7180 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.7028 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6480 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      1.7728 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6704 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9587 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8766 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.5600 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4410 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8118 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5400 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END Q
    PIN D
        AntennaGateArea              0.1872 ;
        AntennaPartialMetalArea      0.7049 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6228 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.7135 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6390 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFSRXL
MACRO SDFFSRX4
    PIN SN
        AntennaGateArea              0.9792 ;
        AntennaPartialMetalArea      4.3586 LAYER met1 ;
        AntennaPartialMetalSideArea  3.6000 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.7957 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6912 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.3024 ;
        AntennaPartialMetalArea      1.6308 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5300 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.4644 ;
        AntennaPartialMetalArea      0.6057 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5076 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.8800 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4500 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.7880 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4086 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END Q
    PIN D
        AntennaGateArea              0.1872 ;
        AntennaPartialMetalArea      0.6530 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6084 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.3060 ;
        AntennaPartialMetalArea      0.6206 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5814 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFSRX4
MACRO SDFFSRX2
    PIN SN
        AntennaGateArea              0.5328 ;
        AntennaPartialMetalArea      3.1596 LAYER met1 ;
        AntennaPartialMetalSideArea  2.5740 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7791 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6912 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      1.6769 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6362 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.8260 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7200 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.5976 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4698 LAYER met1 ;
        AntennaDiffArea              1.4700 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.9836 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6660 LAYER met1 ;
        AntennaDiffArea              1.4700 ;
    END Q
    PIN D
        AntennaGateArea              0.1188 ;
        AntennaPartialMetalArea      0.6912 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6030 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.8298 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6606 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFSRX2
MACRO SDFFSRX1
    PIN SN
        AntennaGateArea              0.3312 ;
        AntennaPartialMetalArea      3.2393 LAYER met1 ;
        AntennaPartialMetalSideArea  2.6514 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7783 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6912 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2376 ;
        AntennaPartialMetalArea      1.6827 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6434 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.8313 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7326 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.1684 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8964 LAYER met1 ;
        AntennaDiffArea              0.7743 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8179 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5958 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN D
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      0.6846 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6066 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.7181 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6174 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFSRX1
MACRO SDFFSHQXL
    PIN SN
        AntennaGateArea              0.5112 ;
        AntennaPartialMetalArea      4.3825 LAYER met1 ;
        AntennaPartialMetalSideArea  3.4038 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9013 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8334 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.3024 ;
        AntennaPartialMetalArea      1.9430 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8702 LAYER met1 ;
    END SE
    PIN Q
        AntennaPartialMetalArea      0.9094 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6912 LAYER met1 ;
        AntennaDiffArea              0.6624 ;
    END Q
    PIN D
        AntennaGateArea              0.2016 ;
        AntennaPartialMetalArea      0.6740 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5868 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.6211 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5598 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFSHQXL
MACRO SDFFSHQX4
    PIN SN
        AntennaGateArea              1.7028 ;
        AntennaPartialMetalArea      6.3668 LAYER met1 ;
        AntennaPartialMetalSideArea  4.5972 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      1.1128 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9450 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.3204 ;
        AntennaPartialMetalArea      1.8757 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7946 LAYER met1 ;
    END SE
    PIN Q
        AntennaPartialMetalArea      3.0493 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8072 LAYER met1 ;
        AntennaDiffArea              3.2540 ;
    END Q
    PIN D
        AntennaGateArea              0.2304 ;
        AntennaPartialMetalArea      0.7034 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5994 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.4428 ;
        AntennaPartialMetalArea      0.5874 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5436 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFSHQX4
MACRO SDFFSHQX2
    PIN SN
        AntennaGateArea              0.9630 ;
        AntennaPartialMetalArea      4.6641 LAYER met1 ;
        AntennaPartialMetalSideArea  3.7458 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8139 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7146 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2664 ;
        AntennaPartialMetalArea      1.7567 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6542 LAYER met1 ;
    END SE
    PIN Q
        AntennaPartialMetalArea      0.8516 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5616 LAYER met1 ;
        AntennaDiffArea              1.4889 ;
    END Q
    PIN D
        AntennaGateArea              0.1404 ;
        AntennaPartialMetalArea      0.7829 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6876 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.6648 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5868 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFSHQX2
MACRO SDFFSHQX1
    PIN SN
        AntennaGateArea              0.5688 ;
        AntennaPartialMetalArea      4.1157 LAYER met1 ;
        AntennaPartialMetalSideArea  3.1932 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      1.1459 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9738 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2376 ;
        AntennaPartialMetalArea      1.9430 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8702 LAYER met1 ;
    END SE
    PIN Q
        AntennaPartialMetalArea      0.9765 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7110 LAYER met1 ;
        AntennaDiffArea              0.9380 ;
    END Q
    PIN D
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      0.7859 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6768 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2016 ;
        AntennaPartialMetalArea      0.6256 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5778 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFSHQX1
MACRO SDFFSXL
    PIN SN
        AntennaGateArea              0.2808 ;
        AntennaPartialMetalArea      2.4372 LAYER met1 ;
        AntennaPartialMetalSideArea  2.3328 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9309 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8100 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.3024 ;
        AntennaPartialMetalArea      1.7385 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6380 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      1.3153 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9666 LAYER met1 ;
        AntennaDiffArea              0.5874 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.7070 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4752 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END Q
    PIN D
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.8215 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6948 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.5980 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5328 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFSXL
MACRO SDFFSX4
    PIN SN
        AntennaGateArea              0.9288 ;
        AntennaPartialMetalArea      3.1887 LAYER met1 ;
        AntennaPartialMetalSideArea  3.1230 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9075 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7650 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2592 ;
        AntennaPartialMetalArea      1.8316 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7100 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      1.1518 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4644 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.2643 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5040 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END Q
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8001 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7236 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.6103 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5166 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFSX4
MACRO SDFFSX2
    PIN SN
        AntennaGateArea              0.5220 ;
        AntennaPartialMetalArea      2.3357 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2752 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9286 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8046 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2376 ;
        AntennaPartialMetalArea      1.8020 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7316 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      0.8237 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5706 LAYER met1 ;
        AntennaDiffArea              1.3927 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.3050 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8136 LAYER met1 ;
        AntennaDiffArea              1.5480 ;
    END Q
    PIN D
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      0.8170 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7380 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.6670 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5616 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFSX2
MACRO SDFFSX1
    PIN SN
        AntennaGateArea              0.3348 ;
        AntennaPartialMetalArea      2.3837 LAYER met1 ;
        AntennaPartialMetalSideArea  2.3220 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9194 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8100 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2376 ;
        AntennaPartialMetalArea      1.7316 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6650 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      1.4336 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0476 LAYER met1 ;
        AntennaDiffArea              0.7732 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6460 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4716 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN D
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      0.8528 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7344 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.7145 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6120 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFSX1
MACRO SDFFRHQXL
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9742 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8550 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.3024 ;
        AntennaPartialMetalArea      1.6910 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6236 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.1260 ;
        AntennaPartialMetalArea      0.9604 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8586 LAYER met1 ;
    END RN
    PIN Q
        AntennaPartialMetalArea      1.0446 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7506 LAYER met1 ;
        AntennaDiffArea              0.8483 ;
    END Q
    PIN D
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.7220 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6444 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6320 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5472 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFRHQXL
MACRO SDFFRHQX4
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9202 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8334 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.3384 ;
        AntennaPartialMetalArea      1.8996 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6074 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.7380 ;
        AntennaPartialMetalArea      1.0394 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9342 LAYER met1 ;
    END RN
    PIN Q
        AntennaPartialMetalArea      3.0205 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6902 LAYER met1 ;
        AntennaDiffArea              2.8368 ;
    END Q
    PIN D
        AntennaGateArea              0.2628 ;
        AntennaPartialMetalArea      0.8767 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7920 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.4788 ;
        AntennaPartialMetalArea      0.6908 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5598 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFRHQX4
MACRO SDFFRHQX2
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9423 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8910 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      1.6898 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6056 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.4140 ;
        AntennaPartialMetalArea      0.6760 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5940 LAYER met1 ;
    END RN
    PIN Q
        AntennaPartialMetalArea      1.2132 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8316 LAYER met1 ;
        AntennaDiffArea              1.4040 ;
    END Q
    PIN D
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.7614 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6750 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2988 ;
        AntennaPartialMetalArea      0.5606 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4842 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFRHQX2
MACRO SDFFRHQX1
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9423 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8910 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      1.7186 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6344 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.2628 ;
        AntennaPartialMetalArea      0.8268 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7398 LAYER met1 ;
    END RN
    PIN Q
        AntennaPartialMetalArea      1.2210 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8802 LAYER met1 ;
        AntennaDiffArea              0.9720 ;
    END Q
    PIN D
        AntennaGateArea              0.1188 ;
        AntennaPartialMetalArea      0.7614 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6750 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2052 ;
        AntennaPartialMetalArea      0.5840 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5076 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFRHQX1
MACRO SDFFRXL
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9817 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8640 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.3024 ;
        AntennaPartialMetalArea      1.7576 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6668 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6449 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5850 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.2640 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9324 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.5979 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4536 LAYER met1 ;
        AntennaDiffArea              0.6339 ;
    END Q
    PIN D
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.8348 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7506 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1260 ;
        AntennaPartialMetalArea      0.9018 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8046 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFRXL
MACRO SDFFRX4
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8012 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6894 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      1.5842 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5246 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.4068 ;
        AntennaPartialMetalArea      1.0354 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9000 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.9546 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4752 LAYER met1 ;
        AntennaDiffArea              1.4157 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8764 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4392 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END Q
    PIN D
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.9539 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8568 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.5831 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5058 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFRX4
MACRO SDFFRX2
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9174 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8298 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2412 ;
        AntennaPartialMetalArea      1.6744 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6110 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      0.7620 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5832 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.9294 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5994 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.1627 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7164 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Q
    PIN D
        AntennaGateArea              0.1116 ;
        AntennaPartialMetalArea      0.9191 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7920 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.6544 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5472 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFRX2
MACRO SDFFRX1
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9925 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8748 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2412 ;
        AntennaPartialMetalArea      1.8388 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7424 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.6683 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5922 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.3015 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9594 LAYER met1 ;
        AntennaDiffArea              0.7776 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6457 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4716 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN D
        AntennaGateArea              0.1116 ;
        AntennaPartialMetalArea      0.8862 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7884 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.7362 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6390 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFRX1
MACRO SDFFNSRXL
    PIN SN
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      3.3774 LAYER met1 ;
        AntennaPartialMetalSideArea  2.7288 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.7160 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6606 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      1.7638 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6614 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9639 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8802 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.7811 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6084 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6124 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4554 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END Q
    PIN D
        AntennaGateArea              0.1872 ;
        AntennaPartialMetalArea      0.7049 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6228 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.6560 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6156 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END SDFFNSRXL
MACRO SDFFNSRX4
    PIN SN
        AntennaGateArea              0.9792 ;
        AntennaPartialMetalArea      4.2695 LAYER met1 ;
        AntennaPartialMetalSideArea  3.5208 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.7551 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6966 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2988 ;
        AntennaPartialMetalArea      1.6273 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5210 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.4572 ;
        AntennaPartialMetalArea      0.7511 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6498 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.9236 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4266 LAYER met1 ;
        AntennaDiffArea              1.4232 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.2160 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4662 LAYER met1 ;
        AntennaDiffArea              1.4232 ;
    END Q
    PIN D
        AntennaGateArea              0.1872 ;
        AntennaPartialMetalArea      0.6520 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6084 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.3060 ;
        AntennaPartialMetalArea      0.6827 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5742 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END SDFFNSRX4
MACRO SDFFNSRX2
    PIN SN
        AntennaGateArea              0.5328 ;
        AntennaPartialMetalArea      3.1839 LAYER met1 ;
        AntennaPartialMetalSideArea  2.6064 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8364 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7362 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      1.6719 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6326 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.8444 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7254 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.7232 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5040 LAYER met1 ;
        AntennaDiffArea              1.7157 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.2744 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7776 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Q
    PIN D
        AntennaGateArea              0.1188 ;
        AntennaPartialMetalArea      0.7018 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6084 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.6566 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6048 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END SDFFNSRX2
MACRO SDFFNSRX1
    PIN SN
        AntennaGateArea              0.3312 ;
        AntennaPartialMetalArea      3.2276 LAYER met1 ;
        AntennaPartialMetalSideArea  2.6748 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8364 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7362 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2376 ;
        AntennaPartialMetalArea      1.6827 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6434 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.8445 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7308 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.9173 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7308 LAYER met1 ;
        AntennaDiffArea              0.7740 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6480 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4734 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN D
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      0.7616 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6372 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.6638 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6120 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END SDFFNSRX1
MACRO SDFFNSXL
    PIN SN
        AntennaGateArea              0.2808 ;
        AntennaPartialMetalArea      2.4945 LAYER met1 ;
        AntennaPartialMetalSideArea  2.3904 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9521 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8172 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.3024 ;
        AntennaPartialMetalArea      1.7457 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6452 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      1.3153 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9666 LAYER met1 ;
        AntennaDiffArea              0.5874 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6870 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4662 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END Q
    PIN D
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.8037 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6858 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6286 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5634 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END SDFFNSXL
MACRO SDFFNSX4
    PIN SN
        AntennaGateArea              0.9288 ;
        AntennaPartialMetalArea      3.3061 LAYER met1 ;
        AntennaPartialMetalSideArea  3.2274 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9103 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7866 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2592 ;
        AntennaPartialMetalArea      1.8511 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7442 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      1.3078 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6336 LAYER met1 ;
        AntennaDiffArea              1.5681 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.0182 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5292 LAYER met1 ;
        AntennaDiffArea              1.5681 ;
    END Q
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8056 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7254 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.5807 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5040 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END SDFFNSX4
MACRO SDFFNSX2
    PIN SN
        AntennaGateArea              0.5220 ;
        AntennaPartialMetalArea      2.4218 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2932 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9404 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7956 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2376 ;
        AntennaPartialMetalArea      1.9242 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7640 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      0.8119 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5652 LAYER met1 ;
        AntennaDiffArea              1.4064 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.2902 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8136 LAYER met1 ;
        AntennaDiffArea              1.5480 ;
    END Q
    PIN D
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      0.7763 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6930 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.6579 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5436 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END SDFFNSX2
MACRO SDFFNSX1
    PIN SN
        AntennaGateArea              0.3348 ;
        AntennaPartialMetalArea      2.4003 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2734 LAYER met1 ;
    END SN
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9056 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8298 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2376 ;
        AntennaPartialMetalArea      1.7779 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6884 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      1.3524 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9972 LAYER met1 ;
        AntennaDiffArea              0.7687 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8116 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4446 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN D
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      0.8896 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7704 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.5944 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5292 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END SDFFNSX1
MACRO SDFFNRXL
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9992 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8766 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.3024 ;
        AntennaPartialMetalArea      1.7121 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6182 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7918 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6894 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.2774 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9630 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.5361 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4320 LAYER met1 ;
        AntennaDiffArea              0.6699 ;
    END Q
    PIN D
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.8628 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7650 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1260 ;
        AntennaPartialMetalArea      0.5992 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5364 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END SDFFNRXL
MACRO SDFFNRX4
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      1.0052 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8982 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      1.8176 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7370 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.3960 ;
        AntennaPartialMetalArea      1.0554 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9486 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.9744 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4806 LAYER met1 ;
        AntennaDiffArea              1.6362 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.0082 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5058 LAYER met1 ;
        AntennaDiffArea              1.6362 ;
    END Q
    PIN D
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.8276 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7452 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.6065 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5292 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END SDFFNRX4
MACRO SDFFNRX2
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9174 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8298 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2412 ;
        AntennaPartialMetalArea      1.6692 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6110 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      0.7620 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5832 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.9294 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5994 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.1594 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7164 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Q
    PIN D
        AntennaGateArea              0.1116 ;
        AntennaPartialMetalArea      0.9191 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7920 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.6544 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5472 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END SDFFNRX2
MACRO SDFFNRX1
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      1.0258 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9072 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2412 ;
        AntennaPartialMetalArea      1.7670 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6992 LAYER met1 ;
    END SE
    PIN RN
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.7846 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6822 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.3099 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9828 LAYER met1 ;
        AntennaDiffArea              0.7776 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.5841 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4662 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN D
        AntennaGateArea              0.1116 ;
        AntennaPartialMetalArea      0.9657 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8442 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.6561 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6084 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END SDFFNRX1
MACRO SDFFNXL
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      1.2791 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0710 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.3024 ;
        AntennaPartialMetalArea      1.8605 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4544 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      0.6432 LAYER met1 ;
        AntennaPartialMetalSideArea  0.3978 LAYER met1 ;
        AntennaDiffArea              0.6564 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.1028 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8280 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END Q
    PIN D
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.8756 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7614 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6169 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5292 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END SDFFNXL
MACRO SDFFNX4
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9918 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8748 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.3312 ;
        AntennaPartialMetalArea      2.0005 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6596 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      0.8080 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4176 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8760 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4482 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END Q
    PIN D
        AntennaGateArea              0.2340 ;
        AntennaPartialMetalArea      0.8554 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7434 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.4788 ;
        AntennaPartialMetalArea      0.7582 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5976 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END SDFFNX4
MACRO SDFFNX2
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      1.2608 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0638 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2592 ;
        AntennaPartialMetalArea      1.8229 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4400 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      1.0742 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7146 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.1225 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8442 LAYER met1 ;
        AntennaDiffArea              1.0500 ;
    END Q
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7903 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7254 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.6081 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5256 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END SDFFNX2
MACRO SDFFNX1
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      1.2661 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0674 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2376 ;
        AntennaPartialMetalArea      1.8310 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4418 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      0.8220 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4500 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.2313 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9054 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN D
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      0.8417 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7398 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.5784 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5148 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END SDFFNX1
MACRO SDFFHQXL
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9870 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8892 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2808 ;
        AntennaPartialMetalArea      1.8252 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7586 LAYER met1 ;
    END SE
    PIN Q
        AntennaPartialMetalArea      1.0804 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8496 LAYER met1 ;
        AntennaDiffArea              0.6853 ;
    END Q
    PIN D
        AntennaGateArea              0.1764 ;
        AntennaPartialMetalArea      0.7440 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6786 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.6580 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6138 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFHQXL
MACRO SDFFHQX4
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      1.2297 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0944 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2952 ;
        AntennaPartialMetalArea      2.0969 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6812 LAYER met1 ;
    END SE
    PIN Q
        AntennaPartialMetalArea      1.4154 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7308 LAYER met1 ;
        AntennaDiffArea              1.7640 ;
    END Q
    PIN D
        AntennaGateArea              0.1872 ;
        AntennaPartialMetalArea      0.8523 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7650 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.3960 ;
        AntennaPartialMetalArea      0.7016 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6354 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFHQX4
MACRO SDFFHQX2
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9228 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8550 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      1.8527 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7694 LAYER met1 ;
    END SE
    PIN Q
        AntennaPartialMetalArea      0.8566 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6354 LAYER met1 ;
        AntennaDiffArea              1.3252 ;
    END Q
    PIN D
        AntennaGateArea              0.1188 ;
        AntennaPartialMetalArea      0.8151 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7578 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.6380 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5850 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFHQX2
MACRO SDFFHQX1
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9300 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8622 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2376 ;
        AntennaPartialMetalArea      1.8769 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7964 LAYER met1 ;
    END SE
    PIN Q
        AntennaPartialMetalArea      1.1582 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8712 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN D
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      0.8726 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7614 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.6464 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6012 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFHQX1
MACRO SDFFXL
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      1.2850 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0710 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.3024 ;
        AntennaPartialMetalArea      1.9048 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4526 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      0.6432 LAYER met1 ;
        AntennaPartialMetalSideArea  0.3978 LAYER met1 ;
        AntennaDiffArea              0.6564 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.1055 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8244 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END Q
    PIN D
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.8788 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7632 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6169 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5292 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFXL
MACRO SDFFX4
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9918 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8748 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.3276 ;
        AntennaPartialMetalArea      2.0111 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6632 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      1.1647 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5112 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.0687 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4734 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END Q
    PIN D
        AntennaGateArea              0.2340 ;
        AntennaPartialMetalArea      0.8590 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7470 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.4788 ;
        AntennaPartialMetalArea      0.7582 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5976 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFX4
MACRO SDFFX2
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      1.2642 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0620 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2592 ;
        AntennaPartialMetalArea      1.8093 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4400 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      1.0750 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7146 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.2297 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8442 LAYER met1 ;
        AntennaDiffArea              1.0500 ;
    END Q
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7877 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7254 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.6081 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5256 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFX2
MACRO SDFFX1
    PIN SI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      1.2948 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0818 LAYER met1 ;
    END SI
    PIN SE
        AntennaGateArea              0.2376 ;
        AntennaPartialMetalArea      1.8621 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4526 LAYER met1 ;
    END SE
    PIN QN
        AntennaPartialMetalArea      0.7705 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5382 LAYER met1 ;
        AntennaDiffArea              0.7860 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.4354 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9846 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN D
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      0.8717 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7632 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.6169 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5292 LAYER met1 ;
    END CK
    PIN GND
    END GND
END SDFFX1
MACRO RSLATNXL
    PIN SN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6728 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6066 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7712 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7128 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.8090 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5382 LAYER met1 ;
        AntennaDiffArea              0.5628 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8352 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5976 LAYER met1 ;
        AntennaDiffArea              0.5628 ;
    END Q
    PIN GND
    END GND
END RSLATNXL
MACRO RSLATNX4
    PIN SN
        AntennaGateArea              0.3924 ;
        AntennaPartialMetalArea      0.6812 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5580 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.3852 ;
        AntennaPartialMetalArea      0.5818 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5094 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.0344 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4482 LAYER met1 ;
        AntennaDiffArea              1.7871 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8120 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4194 LAYER met1 ;
        AntennaDiffArea              1.4157 ;
    END Q
    PIN GND
    END GND
END RSLATNX4
MACRO RSLATNX2
    PIN SN
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.6290 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5508 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.6363 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5688 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.0954 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7380 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.0073 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6840 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Q
    PIN GND
    END GND
END RSLATNX2
MACRO RSLATNX1
    PIN SN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7016 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6354 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8000 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7416 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.8090 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5382 LAYER met1 ;
        AntennaDiffArea              0.7740 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8352 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5976 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN GND
    END GND
END RSLATNX1
MACRO RSLATXL
    PIN S
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6125 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5328 LAYER met1 ;
    END S
    PIN R
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8146 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7272 LAYER met1 ;
    END R
    PIN QN
        AntennaPartialMetalArea      0.7224 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5238 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.9842 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6732 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END Q
    PIN GND
    END GND
END RSLATXL
MACRO RSLATX4
    PIN S
        AntennaGateArea              0.3492 ;
        AntennaPartialMetalArea      0.7016 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6048 LAYER met1 ;
    END S
    PIN R
        AntennaGateArea              0.3492 ;
        AntennaPartialMetalArea      0.6342 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5400 LAYER met1 ;
    END R
    PIN QN
        AntennaPartialMetalArea      0.8598 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4374 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.2321 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6336 LAYER met1 ;
        AntennaDiffArea              1.4292 ;
    END Q
    PIN GND
    END GND
END RSLATX4
MACRO RSLATX2
    PIN S
        AntennaGateArea              0.1692 ;
        AntennaPartialMetalArea      0.5885 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5112 LAYER met1 ;
    END S
    PIN R
        AntennaGateArea              0.1692 ;
        AntennaPartialMetalArea      0.7586 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6678 LAYER met1 ;
    END R
    PIN QN
        AntennaPartialMetalArea      1.0722 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7038 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.9169 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6786 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Q
    PIN GND
    END GND
END RSLATX2
MACRO RSLATX1
    PIN S
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6010 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5166 LAYER met1 ;
    END S
    PIN R
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8300 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7200 LAYER met1 ;
    END R
    PIN QN
        AntennaPartialMetalArea      0.8068 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5886 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8650 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6030 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN GND
    END GND
END RSLATX1
MACRO OR4XL
    PIN Y
        AntennaPartialMetalArea      0.8540 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6138 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END Y
    PIN D
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.8200 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6534 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.6829 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6012 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.7314 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6696 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.7989 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7092 LAYER met1 ;
    END A
    PIN GND
    END GND
END OR4XL
MACRO OR4X4
    PIN Y
        AntennaPartialMetalArea      0.8134 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4158 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END Y
    PIN D
        AntennaGateArea              0.6408 ;
        AntennaPartialMetalArea      2.4494 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9926 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.6408 ;
        AntennaPartialMetalArea      2.2384 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7784 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.6408 ;
        AntennaPartialMetalArea      1.5232 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2546 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.6408 ;
        AntennaPartialMetalArea      1.0226 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8712 LAYER met1 ;
    END A
    PIN GND
    END GND
END OR4X4
MACRO OR4X2
    PIN Y
        AntennaPartialMetalArea      1.3431 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7758 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Y
    PIN D
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      0.7146 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6156 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      0.6568 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5760 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      0.6794 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6264 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      0.7896 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6948 LAYER met1 ;
    END A
    PIN GND
    END GND
END OR4X2
MACRO OR4X1
    PIN Y
        AntennaPartialMetalArea      0.8732 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6138 LAYER met1 ;
        AntennaDiffArea              0.7740 ;
    END Y
    PIN D
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.8112 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6498 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.6826 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5994 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.6974 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6444 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.7873 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7056 LAYER met1 ;
    END A
    PIN GND
    END GND
END OR4X1
MACRO OR3XL
    PIN Y
        AntennaPartialMetalArea      0.7684 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5580 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END Y
    PIN C
        AntennaGateArea              0.1728 ;
        AntennaPartialMetalArea      0.7832 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6372 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.1728 ;
        AntennaPartialMetalArea      0.7111 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6084 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.1728 ;
        AntennaPartialMetalArea      0.6428 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5832 LAYER met1 ;
    END A
    PIN GND
    END GND
END OR3XL
MACRO OR3X4
    PIN Y
        AntennaPartialMetalArea      0.8645 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4392 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END Y
    PIN C
        AntennaGateArea              0.5760 ;
        AntennaPartialMetalArea      1.8354 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5336 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.5760 ;
        AntennaPartialMetalArea      1.3234 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1448 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5760 ;
        AntennaPartialMetalArea      0.8177 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7398 LAYER met1 ;
    END A
    PIN GND
    END GND
END OR3X4
MACRO OR3X2
    PIN Y
        AntennaPartialMetalArea      1.2626 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7848 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Y
    PIN C
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      0.7290 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6300 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      0.6591 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5904 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      0.6756 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5958 LAYER met1 ;
    END A
    PIN GND
    END GND
END OR3X2
MACRO OR3X1
    PIN Y
        AntennaPartialMetalArea      0.8100 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6120 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Y
    PIN C
        AntennaGateArea              0.1728 ;
        AntennaPartialMetalArea      0.7832 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6372 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.1728 ;
        AntennaPartialMetalArea      0.7064 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6066 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.1728 ;
        AntennaPartialMetalArea      0.6451 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5850 LAYER met1 ;
    END A
    PIN GND
    END GND
END OR3X1
MACRO OR2XL
    PIN Y
        AntennaPartialMetalArea      0.7017 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5130 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END Y
    PIN B
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.7750 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6534 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      1.0080 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8766 LAYER met1 ;
    END A
    PIN GND
    END GND
END OR2XL
MACRO OR2X4
    PIN Y
        AntennaPartialMetalArea      0.8941 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4482 LAYER met1 ;
        AntennaDiffArea              1.4112 ;
    END Y
    PIN B
        AntennaGateArea              0.4968 ;
        AntennaPartialMetalArea      0.6117 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5382 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.4968 ;
        AntennaPartialMetalArea      0.6651 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5634 LAYER met1 ;
    END A
    PIN GND
    END GND
END OR2X4
MACRO OR2X2
    PIN Y
        AntennaPartialMetalArea      0.9897 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7074 LAYER met1 ;
        AntennaDiffArea              1.5960 ;
    END Y
    PIN B
        AntennaGateArea              0.2592 ;
        AntennaPartialMetalArea      0.6956 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5778 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.2592 ;
        AntennaPartialMetalArea      0.6824 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5958 LAYER met1 ;
    END A
    PIN GND
    END GND
END OR2X2
MACRO OR2X1
    PIN Y
        AntennaPartialMetalArea      0.7297 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5310 LAYER met1 ;
        AntennaDiffArea              0.7890 ;
    END Y
    PIN B
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.7750 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6534 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.9954 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8712 LAYER met1 ;
    END A
    PIN GND
    END GND
END OR2X1
MACRO OAI33XL
    PIN Y
        AntennaPartialMetalArea      2.0364 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3914 LAYER met1 ;
        AntennaDiffArea              1.3804 ;
    END Y
    PIN B2
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.8757 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7434 LAYER met1 ;
    END B2
    PIN B1
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.7284 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6552 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.8210 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6912 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.8125 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7200 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.7312 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6264 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.7167 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6354 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI33XL
MACRO OAI33X4
    PIN Y
        AntennaPartialMetalArea      0.9632 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5616 LAYER met1 ;
        AntennaDiffArea              1.7277 ;
    END Y
    PIN B2
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.8574 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7668 LAYER met1 ;
    END B2
    PIN B1
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.7369 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6444 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.7995 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7110 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.7695 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6642 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.7322 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6588 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.8145 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7272 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI33X4
MACRO OAI33X2
    PIN Y
        AntennaPartialMetalArea      2.8997 LAYER met1 ;
        AntennaPartialMetalSideArea  2.1924 LAYER met1 ;
        AntennaDiffArea              3.3005 ;
    END Y
    PIN B2
        AntennaGateArea              0.7938 ;
        AntennaPartialMetalArea      2.1900 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6614 LAYER met1 ;
    END B2
    PIN B1
        AntennaGateArea              0.7938 ;
        AntennaPartialMetalArea      1.3283 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1700 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.7938 ;
        AntennaPartialMetalArea      0.8732 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7938 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.7938 ;
        AntennaPartialMetalArea      2.2717 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8270 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.7938 ;
        AntennaPartialMetalArea      1.3281 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1592 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.7938 ;
        AntennaPartialMetalArea      0.8007 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6966 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI33X2
MACRO OAI33X1
    PIN Y
        AntennaPartialMetalArea      1.8262 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3194 LAYER met1 ;
        AntennaDiffArea              1.7322 ;
    END Y
    PIN B2
        AntennaGateArea              0.3924 ;
        AntennaPartialMetalArea      0.7887 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6588 LAYER met1 ;
    END B2
    PIN B1
        AntennaGateArea              0.3924 ;
        AntennaPartialMetalArea      0.6767 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6012 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.3924 ;
        AntennaPartialMetalArea      0.7472 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6408 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.3924 ;
        AntennaPartialMetalArea      0.7639 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6714 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.3924 ;
        AntennaPartialMetalArea      0.6691 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5778 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.3924 ;
        AntennaPartialMetalArea      0.7260 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5832 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI33X1
MACRO OAI32XL
    PIN Y
        AntennaPartialMetalArea      1.4784 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0800 LAYER met1 ;
        AntennaDiffArea              0.9114 ;
    END Y
    PIN B1
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.8046 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7272 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.8444 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7524 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.8503 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6984 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.7260 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6534 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.8248 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7128 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI32XL
MACRO OAI32X4
    PIN Y
        AntennaPartialMetalArea      1.1272 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5706 LAYER met1 ;
        AntennaDiffArea              1.7277 ;
    END Y
    PIN B1
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      0.7610 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6516 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      0.9185 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7848 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.8467 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7380 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.7089 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6174 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.7254 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6462 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI32X4
MACRO OAI32X2
    PIN Y
        AntennaPartialMetalArea      2.6304 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8684 LAYER met1 ;
        AntennaDiffArea              2.9891 ;
    END Y
    PIN B1
        AntennaGateArea              0.7218 ;
        AntennaPartialMetalArea      1.4507 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2150 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.7218 ;
        AntennaPartialMetalArea      0.7985 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7416 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.7938 ;
        AntennaPartialMetalArea      2.1852 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6470 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.7938 ;
        AntennaPartialMetalArea      1.3175 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1592 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.7938 ;
        AntennaPartialMetalArea      0.8704 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7938 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI32X2
MACRO OAI32X1
    PIN Y
        AntennaPartialMetalArea      1.3484 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0350 LAYER met1 ;
        AntennaDiffArea              1.2760 ;
    END Y
    PIN B1
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7560 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6876 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.8330 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6822 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.3960 ;
        AntennaPartialMetalArea      0.7996 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6588 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.3960 ;
        AntennaPartialMetalArea      0.6856 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6138 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.3960 ;
        AntennaPartialMetalArea      0.7852 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6732 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI32X1
MACRO OAI31XL
    PIN Y
        AntennaPartialMetalArea      1.0746 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7776 LAYER met1 ;
        AntennaDiffArea              0.9368 ;
    END Y
    PIN B0
        AntennaGateArea              0.2160 ;
        AntennaPartialMetalArea      0.7372 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6210 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.7420 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6084 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.6161 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5742 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.8592 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7578 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI31XL
MACRO OAI31X4
    PIN Y
        AntennaPartialMetalArea      1.0278 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5778 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END Y
    PIN B0
        AntennaGateArea              0.1944 ;
        AntennaPartialMetalArea      0.8690 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7920 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.8519 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7272 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.7089 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6174 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.7680 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6588 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI31X4
MACRO OAI31X2
    PIN Y
        AntennaPartialMetalArea      1.5441 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1466 LAYER met1 ;
        AntennaDiffArea              1.7820 ;
    END Y
    PIN B0
        AntennaGateArea              0.6120 ;
        AntennaPartialMetalArea      1.2452 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0134 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.8100 ;
        AntennaPartialMetalArea      2.1964 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8630 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.8100 ;
        AntennaPartialMetalArea      1.5744 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3518 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.8100 ;
        AntennaPartialMetalArea      1.0558 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9072 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI31X2
MACRO OAI31X1
    PIN Y
        AntennaPartialMetalArea      1.0502 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7578 LAYER met1 ;
        AntennaDiffArea              1.2320 ;
    END Y
    PIN B0
        AntennaGateArea              0.3060 ;
        AntennaPartialMetalArea      0.6654 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6138 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.3960 ;
        AntennaPartialMetalArea      0.7472 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6066 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.3960 ;
        AntennaPartialMetalArea      0.6298 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5760 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.3960 ;
        AntennaPartialMetalArea      0.8496 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7488 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI31X1
MACRO OAI2BB2XL
    PIN Y
        AntennaPartialMetalArea      1.2340 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9072 LAYER met1 ;
        AntennaDiffArea              0.7228 ;
    END Y
    PIN B1
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7779 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7038 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.8242 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7524 LAYER met1 ;
    END B0
    PIN A1N
        AntennaGateArea              0.1404 ;
        AntennaPartialMetalArea      0.6495 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5778 LAYER met1 ;
    END A1N
    PIN A0N
        AntennaGateArea              0.1404 ;
        AntennaPartialMetalArea      0.9032 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8172 LAYER met1 ;
    END A0N
    PIN GND
    END GND
END OAI2BB2XL
MACRO OAI2BB2X4
    PIN Y
        AntennaPartialMetalArea      3.5633 LAYER met1 ;
        AntennaPartialMetalSideArea  2.4210 LAYER met1 ;
        AntennaDiffArea              3.8009 ;
    END Y
    PIN B1
        AntennaGateArea              1.4364 ;
        AntennaPartialMetalArea      2.5887 LAYER met1 ;
        AntennaPartialMetalSideArea  2.0700 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              1.4364 ;
        AntennaPartialMetalArea      2.5807 LAYER met1 ;
        AntennaPartialMetalSideArea  2.1942 LAYER met1 ;
    END B0
    PIN A1N
        AntennaGateArea              0.5544 ;
        AntennaPartialMetalArea      1.1082 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9216 LAYER met1 ;
    END A1N
    PIN A0N
        AntennaGateArea              0.5544 ;
        AntennaPartialMetalArea      2.4616 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9566 LAYER met1 ;
    END A0N
    PIN GND
    END GND
END OAI2BB2X4
MACRO OAI2BB2X2
    PIN Y
        AntennaPartialMetalArea      2.0961 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5246 LAYER met1 ;
        AntennaDiffArea              1.8728 ;
    END Y
    PIN B1
        AntennaGateArea              0.7164 ;
        AntennaPartialMetalArea      2.1382 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7586 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.7164 ;
        AntennaPartialMetalArea      1.6786 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6092 LAYER met1 ;
    END B0
    PIN A1N
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.7774 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7074 LAYER met1 ;
    END A1N
    PIN A0N
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.8678 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7182 LAYER met1 ;
    END A0N
    PIN GND
    END GND
END OAI2BB2X2
MACRO OAI2BB2X1
    PIN Y
        AntennaPartialMetalArea      1.1860 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8856 LAYER met1 ;
        AntennaDiffArea              1.0220 ;
    END Y
    PIN B1
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.8210 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6840 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.8092 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7074 LAYER met1 ;
    END B0
    PIN A1N
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.6832 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6084 LAYER met1 ;
    END A1N
    PIN A0N
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      1.0764 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9198 LAYER met1 ;
    END A0N
    PIN GND
    END GND
END OAI2BB2X1
MACRO OAI2BB1XL
    PIN Y
        AntennaPartialMetalArea      0.9508 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7560 LAYER met1 ;
        AntennaDiffArea              0.6624 ;
    END Y
    PIN B0
        AntennaGateArea              0.2160 ;
        AntennaPartialMetalArea      0.8068 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7200 LAYER met1 ;
    END B0
    PIN A1N
        AntennaGateArea              0.1404 ;
        AntennaPartialMetalArea      0.9977 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9360 LAYER met1 ;
    END A1N
    PIN A0N
        AntennaGateArea              0.1404 ;
        AntennaPartialMetalArea      0.7901 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7020 LAYER met1 ;
    END A0N
    PIN GND
    END GND
END OAI2BB1XL
MACRO OAI2BB1X4
    PIN Y
        AntennaPartialMetalArea      2.6925 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2078 LAYER met1 ;
        AntennaDiffArea              2.9522 ;
    END Y
    PIN B0
        AntennaGateArea              1.2348 ;
        AntennaPartialMetalArea      2.2519 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6362 LAYER met1 ;
    END B0
    PIN A1N
        AntennaGateArea              0.5616 ;
        AntennaPartialMetalArea      0.6731 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5850 LAYER met1 ;
    END A1N
    PIN A0N
        AntennaGateArea              0.5616 ;
        AntennaPartialMetalArea      0.7096 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6354 LAYER met1 ;
    END A0N
    PIN GND
    END GND
END OAI2BB1X4
MACRO OAI2BB1X2
    PIN Y
        AntennaPartialMetalArea      1.0243 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6750 LAYER met1 ;
        AntennaDiffArea              1.6586 ;
    END Y
    PIN B0
        AntennaGateArea              0.6192 ;
        AntennaPartialMetalArea      1.3001 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2492 LAYER met1 ;
    END B0
    PIN A1N
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.8432 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6696 LAYER met1 ;
    END A1N
    PIN A0N
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.7803 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6714 LAYER met1 ;
    END A0N
    PIN GND
    END GND
END OAI2BB1X2
MACRO OAI2BB1X1
    PIN Y
        AntennaPartialMetalArea      1.0431 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7560 LAYER met1 ;
        AntennaDiffArea              0.9380 ;
    END Y
    PIN B0
        AntennaGateArea              0.3060 ;
        AntennaPartialMetalArea      0.8222 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6984 LAYER met1 ;
    END B0
    PIN A1N
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      1.0200 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9414 LAYER met1 ;
    END A1N
    PIN A0N
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.7610 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6750 LAYER met1 ;
    END A0N
    PIN GND
    END GND
END OAI2BB1X1
MACRO OAI22XL
    PIN Y
        AntennaPartialMetalArea      1.3820 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0602 LAYER met1 ;
        AntennaDiffArea              0.8120 ;
    END Y
    PIN B1
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7594 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6282 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.8152 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7020 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7860 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6336 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.8550 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7236 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI22XL
MACRO OAI22X4
    PIN Y
        AntennaPartialMetalArea      5.7393 LAYER met1 ;
        AntennaPartialMetalSideArea  3.1464 LAYER met1 ;
        AntennaDiffArea              5.0202 ;
    END Y
    PIN B1
        AntennaGateArea              1.4472 ;
        AntennaPartialMetalArea      1.9107 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6560 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              1.4472 ;
        AntennaPartialMetalArea      2.0242 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6344 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              1.4472 ;
        AntennaPartialMetalArea      2.2353 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7046 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              1.4472 ;
        AntennaPartialMetalArea      2.0143 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6632 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI22X4
MACRO OAI22X2
    PIN Y
        AntennaPartialMetalArea      3.4790 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2914 LAYER met1 ;
        AntennaDiffArea              2.8828 ;
    END Y
    PIN B1
        AntennaGateArea              0.7128 ;
        AntennaPartialMetalArea      1.3750 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9684 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.7128 ;
        AntennaPartialMetalArea      1.8245 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4778 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.7128 ;
        AntennaPartialMetalArea      1.2086 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0494 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.7128 ;
        AntennaPartialMetalArea      1.7949 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4760 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI22X2
MACRO OAI22X1
    PIN Y
        AntennaPartialMetalArea      1.3744 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0440 LAYER met1 ;
        AntennaDiffArea              1.1600 ;
    END Y
    PIN B1
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7712 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6336 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.8120 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7128 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7918 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6282 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.8516 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7110 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI22X1
MACRO OAI222XL
    PIN Y
        AntennaPartialMetalArea      1.9977 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4400 LAYER met1 ;
        AntennaDiffArea              1.3068 ;
    END Y
    PIN C1
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.8813 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7380 LAYER met1 ;
    END C1
    PIN C0
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.8938 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7848 LAYER met1 ;
    END C0
    PIN B1
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.8751 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7326 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.7733 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6588 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.8050 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7254 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.8952 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7650 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI222XL
MACRO OAI222X4
    PIN Y
        AntennaPartialMetalArea      1.1579 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5724 LAYER met1 ;
        AntennaDiffArea              1.7400 ;
    END Y
    PIN C1
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.7534 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6786 LAYER met1 ;
    END C1
    PIN C0
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.7341 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6606 LAYER met1 ;
    END C0
    PIN B1
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.9274 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7722 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.8882 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7218 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.7904 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7020 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.7925 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7236 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI222X4
MACRO OAI222X2
    PIN Y
        AntennaPartialMetalArea      3.4940 LAYER met1 ;
        AntennaPartialMetalSideArea  2.4858 LAYER met1 ;
        AntennaDiffArea              3.1488 ;
    END Y
    PIN C1
        AntennaGateArea              0.7776 ;
        AntennaPartialMetalArea      1.7852 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4724 LAYER met1 ;
    END C1
    PIN C0
        AntennaGateArea              0.7776 ;
        AntennaPartialMetalArea      1.2740 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9702 LAYER met1 ;
    END C0
    PIN B1
        AntennaGateArea              0.7740 ;
        AntennaPartialMetalArea      1.6854 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3662 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.7740 ;
        AntennaPartialMetalArea      1.0979 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8676 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.7956 ;
        AntennaPartialMetalArea      1.8391 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4670 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.7956 ;
        AntennaPartialMetalArea      0.9654 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8028 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI222X2
MACRO OAI222X1
    PIN Y
        AntennaPartialMetalArea      1.8355 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3302 LAYER met1 ;
        AntennaDiffArea              1.8768 ;
    END Y
    PIN C1
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.6484 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5796 LAYER met1 ;
    END C1
    PIN C0
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.8298 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6660 LAYER met1 ;
    END C0
    PIN B1
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.8572 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7002 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.9064 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7974 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.8032 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6642 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.6335 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5436 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI222X1
MACRO OAI221XL
    PIN Y
        AntennaPartialMetalArea      1.6641 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1772 LAYER met1 ;
        AntennaDiffArea              1.1632 ;
    END Y
    PIN C0
        AntennaGateArea              0.2340 ;
        AntennaPartialMetalArea      0.8670 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7560 LAYER met1 ;
    END C0
    PIN B1
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.8827 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6912 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.8488 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6966 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.8981 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7848 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.8469 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7488 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI221XL
MACRO OAI221X4
    PIN Y
        AntennaPartialMetalArea      1.3808 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6642 LAYER met1 ;
        AntennaDiffArea              1.7400 ;
    END Y
    PIN C0
        AntennaGateArea              0.2160 ;
        AntennaPartialMetalArea      0.9510 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8172 LAYER met1 ;
    END C0
    PIN B1
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.8015 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6930 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.8119 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6912 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.9174 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8280 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.8920 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7182 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI221X4
MACRO OAI221X2
    PIN Y
        AntennaPartialMetalArea      2.3118 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6452 LAYER met1 ;
        AntennaDiffArea              2.4324 ;
    END Y
    PIN C0
        AntennaGateArea              0.6696 ;
        AntennaPartialMetalArea      1.1424 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9414 LAYER met1 ;
    END C0
    PIN B1
        AntennaGateArea              0.7776 ;
        AntennaPartialMetalArea      1.7971 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5444 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.7776 ;
        AntennaPartialMetalArea      1.1494 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0062 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.7794 ;
        AntennaPartialMetalArea      1.5138 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2276 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.7794 ;
        AntennaPartialMetalArea      0.8589 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7128 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI221X2
MACRO OAI221X1
    PIN Y
        AntennaPartialMetalArea      1.6859 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1736 LAYER met1 ;
        AntennaDiffArea              1.7472 ;
    END Y
    PIN C0
        AntennaGateArea              0.3348 ;
        AntennaPartialMetalArea      0.6973 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5886 LAYER met1 ;
    END C0
    PIN B1
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.7707 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6570 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.8310 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6768 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.9054 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8118 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.8656 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7632 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI221X1
MACRO OAI21XL
    PIN Y
        AntennaPartialMetalArea      1.0506 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7812 LAYER met1 ;
        AntennaDiffArea              0.7408 ;
    END Y
    PIN B0
        AntennaGateArea              0.2160 ;
        AntennaPartialMetalArea      0.7494 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6642 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7330 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5940 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.6989 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6066 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI21XL
MACRO OAI21X4
    PIN Y
        AntennaPartialMetalArea      3.1083 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2402 LAYER met1 ;
        AntennaDiffArea              3.1612 ;
    END Y
    PIN B0
        AntennaGateArea              1.1808 ;
        AntennaPartialMetalArea      1.2565 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0260 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              1.4580 ;
        AntennaPartialMetalArea      2.3096 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8414 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              1.4580 ;
        AntennaPartialMetalArea      2.3341 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7946 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI21X4
MACRO OAI21X2
    PIN Y
        AntennaPartialMetalArea      1.7801 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2942 LAYER met1 ;
        AntennaDiffArea              1.9460 ;
    END Y
    PIN B0
        AntennaGateArea              0.6084 ;
        AntennaPartialMetalArea      0.8059 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7326 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.7164 ;
        AntennaPartialMetalArea      1.3336 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9936 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.7164 ;
        AntennaPartialMetalArea      1.8467 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4940 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI21X2
MACRO OAI21X1
    PIN Y
        AntennaPartialMetalArea      1.0164 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7308 LAYER met1 ;
        AntennaDiffArea              1.0720 ;
    END Y
    PIN B0
        AntennaGateArea              0.3060 ;
        AntennaPartialMetalArea      0.6088 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5400 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.8410 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6552 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.9352 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7740 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI21X1
MACRO OAI211XL
    PIN Y
        AntennaPartialMetalArea      1.5242 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9990 LAYER met1 ;
        AntennaDiffArea              1.1296 ;
    END Y
    PIN C0
        AntennaGateArea              0.2340 ;
        AntennaPartialMetalArea      0.6238 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5490 LAYER met1 ;
    END C0
    PIN B0
        AntennaGateArea              0.2340 ;
        AntennaPartialMetalArea      0.6532 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5652 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.7909 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6552 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.8912 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7596 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI211XL
MACRO OAI211X4
    PIN Y
        AntennaPartialMetalArea      1.6631 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7704 LAYER met1 ;
        AntennaDiffArea              1.7400 ;
    END Y
    PIN C0
        AntennaGateArea              0.2124 ;
        AntennaPartialMetalArea      0.6596 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5814 LAYER met1 ;
    END C0
    PIN B0
        AntennaGateArea              0.2124 ;
        AntennaPartialMetalArea      0.8886 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8118 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.8422 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7470 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.7196 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6606 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI211X4
MACRO OAI211X2
    PIN Y
        AntennaPartialMetalArea      2.5836 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8882 LAYER met1 ;
        AntennaDiffArea              2.9808 ;
    END Y
    PIN C0
        AntennaGateArea              0.6696 ;
        AntennaPartialMetalArea      1.6578 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3284 LAYER met1 ;
    END C0
    PIN B0
        AntennaGateArea              0.6696 ;
        AntennaPartialMetalArea      0.8233 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7398 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.7740 ;
        AntennaPartialMetalArea      1.3420 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9846 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.7740 ;
        AntennaPartialMetalArea      1.8663 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4796 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI211X2
MACRO OAI211X1
    PIN Y
        AntennaPartialMetalArea      1.4201 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9738 LAYER met1 ;
        AntennaDiffArea              1.6836 ;
    END Y
    PIN C0
        AntennaGateArea              0.3348 ;
        AntennaPartialMetalArea      0.7630 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6588 LAYER met1 ;
    END C0
    PIN B0
        AntennaGateArea              0.3348 ;
        AntennaPartialMetalArea      0.5951 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5256 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.7838 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6282 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.7922 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6876 LAYER met1 ;
    END A0
    PIN GND
    END GND
END OAI211X1
MACRO NOR4BBXL
    PIN Y
        AntennaPartialMetalArea      2.4192 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8018 LAYER met1 ;
        AntennaDiffArea              1.2176 ;
    END Y
    PIN D
        AntennaGateArea              0.2844 ;
        AntennaPartialMetalArea      0.7100 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6570 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.2844 ;
        AntennaPartialMetalArea      0.6644 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5724 LAYER met1 ;
    END C
    PIN BN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6218 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5832 LAYER met1 ;
    END BN
    PIN AN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8902 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7218 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NOR4BBXL
MACRO NOR4BBX4
    PIN Y
        AntennaPartialMetalArea      5.8684 LAYER met1 ;
        AntennaPartialMetalSideArea  4.2570 LAYER met1 ;
        AntennaDiffArea              4.1760 ;
    END Y
    PIN D
        AntennaGateArea              1.4256 ;
        AntennaPartialMetalArea      4.2338 LAYER met1 ;
        AntennaPartialMetalSideArea  3.3534 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              1.4256 ;
        AntennaPartialMetalArea      4.4310 LAYER met1 ;
        AntennaPartialMetalSideArea  3.4992 LAYER met1 ;
    END C
    PIN BN
        AntennaGateArea              0.5832 ;
        AntennaPartialMetalArea      0.6054 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5004 LAYER met1 ;
    END BN
    PIN AN
        AntennaGateArea              0.5832 ;
        AntennaPartialMetalArea      0.6293 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5598 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NOR4BBX4
MACRO NOR4BBX2
    PIN Y
        AntennaPartialMetalArea      3.3150 LAYER met1 ;
        AntennaPartialMetalSideArea  2.4750 LAYER met1 ;
        AntennaDiffArea              2.2712 ;
    END Y
    PIN D
        AntennaGateArea              0.8064 ;
        AntennaPartialMetalArea      2.4106 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9548 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.8064 ;
        AntennaPartialMetalArea      1.8727 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5138 LAYER met1 ;
    END C
    PIN BN
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      0.9273 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8496 LAYER met1 ;
    END BN
    PIN AN
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      0.9104 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6930 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NOR4BBX2
MACRO NOR4BBX1
    PIN Y
        AntennaPartialMetalArea      2.3702 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7946 LAYER met1 ;
        AntennaDiffArea              1.5488 ;
    END Y
    PIN D
        AntennaGateArea              0.4032 ;
        AntennaPartialMetalArea      0.6938 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6408 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.4032 ;
        AntennaPartialMetalArea      0.5992 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5382 LAYER met1 ;
    END C
    PIN BN
        AntennaGateArea              0.1620 ;
        AntennaPartialMetalArea      0.6064 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5652 LAYER met1 ;
    END BN
    PIN AN
        AntennaGateArea              0.1620 ;
        AntennaPartialMetalArea      0.8739 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7074 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NOR4BBX1
MACRO NOR4BXL
    PIN Y
        AntennaPartialMetalArea      1.4108 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0818 LAYER met1 ;
        AntennaDiffArea              1.1686 ;
    END Y
    PIN D
        AntennaGateArea              0.2844 ;
        AntennaPartialMetalArea      0.7691 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6372 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.2844 ;
        AntennaPartialMetalArea      0.6968 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6246 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.2844 ;
        AntennaPartialMetalArea      0.7013 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6228 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8865 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7200 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NOR4BXL
MACRO NOR4BX4
    PIN Y
        AntennaPartialMetalArea      7.5179 LAYER met1 ;
        AntennaPartialMetalSideArea  3.6666 LAYER met1 ;
        AntennaDiffArea              4.1760 ;
    END Y
    PIN D
        AntennaGateArea              1.4256 ;
        AntennaPartialMetalArea      4.2364 LAYER met1 ;
        AntennaPartialMetalSideArea  3.3300 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              1.4256 ;
        AntennaPartialMetalArea      4.3438 LAYER met1 ;
        AntennaPartialMetalSideArea  3.4956 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              1.4256 ;
        AntennaPartialMetalArea      3.7568 LAYER met1 ;
        AntennaPartialMetalSideArea  2.9394 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.5832 ;
        AntennaPartialMetalArea      0.6275 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5580 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NOR4BX4
MACRO NOR4BX2
    PIN Y
        AntennaPartialMetalArea      2.4147 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8234 LAYER met1 ;
        AntennaDiffArea              2.3432 ;
    END Y
    PIN D
        AntennaGateArea              0.8064 ;
        AntennaPartialMetalArea      2.4688 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9134 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.8064 ;
        AntennaPartialMetalArea      1.9008 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5930 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.8064 ;
        AntennaPartialMetalArea      1.4311 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2294 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      0.7585 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6606 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NOR4BX2
MACRO NOR4BX1
    PIN Y
        AntennaPartialMetalArea      1.5746 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1466 LAYER met1 ;
        AntennaDiffArea              1.4432 ;
    END Y
    PIN D
        AntennaGateArea              0.4032 ;
        AntennaPartialMetalArea      0.6920 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6390 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.4032 ;
        AntennaPartialMetalArea      0.5992 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5382 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.4032 ;
        AntennaPartialMetalArea      0.6518 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5796 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.1620 ;
        AntennaPartialMetalArea      0.8919 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7254 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NOR4BX1
MACRO NOR4XL
    PIN Y
        AntennaPartialMetalArea      1.5212 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0872 LAYER met1 ;
        AntennaDiffArea              1.2176 ;
    END Y
    PIN D
        AntennaGateArea              0.2844 ;
        AntennaPartialMetalArea      0.9424 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7020 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.2844 ;
        AntennaPartialMetalArea      0.7220 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6372 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.2844 ;
        AntennaPartialMetalArea      0.6161 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5526 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.2844 ;
        AntennaPartialMetalArea      0.7506 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6426 LAYER met1 ;
    END A
    PIN GND
    END GND
END NOR4XL
MACRO NOR4X4
    PIN Y
        AntennaPartialMetalArea      5.7850 LAYER met1 ;
        AntennaPartialMetalSideArea  3.7782 LAYER met1 ;
        AntennaDiffArea              4.6728 ;
    END Y
    PIN D
        AntennaGateArea              1.4256 ;
        AntennaPartialMetalArea      4.6379 LAYER met1 ;
        AntennaPartialMetalSideArea  3.4488 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              1.4256 ;
        AntennaPartialMetalArea      4.4331 LAYER met1 ;
        AntennaPartialMetalSideArea  3.5496 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              1.4256 ;
        AntennaPartialMetalArea      3.8018 LAYER met1 ;
        AntennaPartialMetalSideArea  2.9430 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              1.4256 ;
        AntennaPartialMetalArea      2.1335 LAYER met1 ;
        AntennaPartialMetalSideArea  2.0610 LAYER met1 ;
    END A
    PIN GND
    END GND
END NOR4X4
MACRO NOR4X2
    PIN Y
        AntennaPartialMetalArea      2.6016 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9584 LAYER met1 ;
        AntennaDiffArea              2.3432 ;
    END Y
    PIN D
        AntennaGateArea              0.8064 ;
        AntennaPartialMetalArea      2.4842 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9170 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.8064 ;
        AntennaPartialMetalArea      1.9401 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6056 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.8064 ;
        AntennaPartialMetalArea      1.4285 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2402 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.8064 ;
        AntennaPartialMetalArea      0.9019 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8118 LAYER met1 ;
    END A
    PIN GND
    END GND
END NOR4X2
MACRO NOR4X1
    PIN Y
        AntennaPartialMetalArea      1.6797 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1466 LAYER met1 ;
        AntennaDiffArea              1.4432 ;
    END Y
    PIN D
        AntennaGateArea              0.4032 ;
        AntennaPartialMetalArea      0.9430 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6840 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.4032 ;
        AntennaPartialMetalArea      0.7316 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6192 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.4032 ;
        AntennaPartialMetalArea      0.6224 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5508 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.4032 ;
        AntennaPartialMetalArea      0.6948 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6120 LAYER met1 ;
    END A
    PIN GND
    END GND
END NOR4X1
MACRO NOR3BXL
    PIN Y
        AntennaPartialMetalArea      1.3258 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9684 LAYER met1 ;
        AntennaDiffArea              1.0606 ;
    END Y
    PIN C
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7652 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6444 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.6673 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5904 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8440 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7254 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NOR3BXL
MACRO NOR3BX4
    PIN Y
        AntennaPartialMetalArea      4.9345 LAYER met1 ;
        AntennaPartialMetalSideArea  2.4192 LAYER met1 ;
        AntennaDiffArea              3.5148 ;
    END Y
    PIN C
        AntennaGateArea              1.2312 ;
        AntennaPartialMetalArea      2.2605 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8594 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              1.2312 ;
        AntennaPartialMetalArea      2.6410 LAYER met1 ;
        AntennaPartialMetalSideArea  2.1024 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.4896 ;
        AntennaPartialMetalArea      0.9998 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8694 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NOR3BX4
MACRO NOR3BX2
    PIN Y
        AntennaPartialMetalArea      2.4156 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4850 LAYER met1 ;
        AntennaDiffArea              2.1560 ;
    END Y
    PIN C
        AntennaGateArea              0.7200 ;
        AntennaPartialMetalArea      2.0724 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7262 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.7200 ;
        AntennaPartialMetalArea      1.4917 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2492 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      0.8053 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6858 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NOR3BX2
MACRO NOR3BX1
    PIN Y
        AntennaPartialMetalArea      1.4613 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0350 LAYER met1 ;
        AntennaDiffArea              1.4120 ;
    END Y
    PIN C
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.6539 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5796 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.6663 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5922 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.1440 ;
        AntennaPartialMetalArea      0.6308 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5598 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NOR3BX1
MACRO NOR3XL
    PIN Y
        AntennaPartialMetalArea      1.6233 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1574 LAYER met1 ;
        AntennaDiffArea              1.0606 ;
    END Y
    PIN C
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.8756 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6570 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.6889 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6228 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7850 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7020 LAYER met1 ;
    END A
    PIN GND
    END GND
END NOR3XL
MACRO NOR3X4
    PIN Y
        AntennaPartialMetalArea      4.6578 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2986 LAYER met1 ;
        AntennaDiffArea              3.4240 ;
    END Y
    PIN C
        AntennaGateArea              1.1880 ;
        AntennaPartialMetalArea      2.8978 LAYER met1 ;
        AntennaPartialMetalSideArea  2.1834 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              1.1880 ;
        AntennaPartialMetalArea      2.6115 LAYER met1 ;
        AntennaPartialMetalSideArea  2.1744 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              1.1880 ;
        AntennaPartialMetalArea      2.3085 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9530 LAYER met1 ;
    END A
    PIN GND
    END GND
END NOR3X4
MACRO NOR3X2
    PIN Y
        AntennaPartialMetalArea      2.5639 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5282 LAYER met1 ;
        AntennaDiffArea              2.5403 ;
    END Y
    PIN C
        AntennaGateArea              0.7200 ;
        AntennaPartialMetalArea      1.7728 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4184 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.7200 ;
        AntennaPartialMetalArea      1.5606 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3140 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.7200 ;
        AntennaPartialMetalArea      0.8524 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7650 LAYER met1 ;
    END A
    PIN GND
    END GND
END NOR3X2
MACRO NOR3X1
    PIN Y
        AntennaPartialMetalArea      1.4698 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0494 LAYER met1 ;
        AntennaDiffArea              1.2872 ;
    END Y
    PIN C
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7917 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6606 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.6851 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6246 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.8044 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7038 LAYER met1 ;
    END A
    PIN GND
    END GND
END NOR3X1
MACRO NOR2BXL
    PIN Y
        AntennaPartialMetalArea      0.8793 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6498 LAYER met1 ;
        AntennaDiffArea              1.0716 ;
    END Y
    PIN B
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      0.7801 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6876 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7384 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6534 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NOR2BXL
MACRO NOR2BX4
    PIN Y
        AntennaPartialMetalArea      3.5022 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7082 LAYER met1 ;
        AntennaDiffArea              2.9274 ;
    END Y
    PIN B
        AntennaGateArea              1.2960 ;
        AntennaPartialMetalArea      1.6543 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4274 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.5148 ;
        AntennaPartialMetalArea      0.7309 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5904 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NOR2BX4
MACRO NOR2BX2
    PIN Y
        AntennaPartialMetalArea      1.5290 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1664 LAYER met1 ;
        AntennaDiffArea              1.4090 ;
    END Y
    PIN B
        AntennaGateArea              0.6480 ;
        AntennaPartialMetalArea      1.5477 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2834 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.2628 ;
        AntennaPartialMetalArea      0.8010 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6606 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NOR2BX2
MACRO NOR2BX1
    PIN Y
        AntennaPartialMetalArea      1.2446 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8658 LAYER met1 ;
        AntennaDiffArea              1.0440 ;
    END Y
    PIN B
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      0.6880 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5994 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6560 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5850 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NOR2BX1
MACRO NOR2XL
    PIN Y
        AntennaPartialMetalArea      1.0691 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7488 LAYER met1 ;
        AntennaDiffArea              0.7344 ;
    END Y
    PIN B
        AntennaGateArea              0.2232 ;
        AntennaPartialMetalArea      0.9646 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6876 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.2232 ;
        AntennaPartialMetalArea      0.7304 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6696 LAYER met1 ;
    END A
    PIN GND
    END GND
END NOR2XL
MACRO NOR2X4
    PIN Y
        AntennaPartialMetalArea      3.5310 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6902 LAYER met1 ;
        AntennaDiffArea              3.1524 ;
    END Y
    PIN B
        AntennaGateArea              1.2960 ;
        AntennaPartialMetalArea      1.7493 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4760 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              1.2960 ;
        AntennaPartialMetalArea      2.0222 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5876 LAYER met1 ;
    END A
    PIN GND
    END GND
END NOR2X4
MACRO NOR2X2
    PIN Y
        AntennaPartialMetalArea      1.6684 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0422 LAYER met1 ;
        AntennaDiffArea              1.9200 ;
    END Y
    PIN B
        AntennaGateArea              0.6480 ;
        AntennaPartialMetalArea      1.4763 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1538 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.6480 ;
        AntennaPartialMetalArea      0.8124 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6858 LAYER met1 ;
    END A
    PIN GND
    END GND
END NOR2X2
MACRO NOR2X1
    PIN Y
        AntennaPartialMetalArea      0.9265 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6732 LAYER met1 ;
        AntennaDiffArea              0.9480 ;
    END Y
    PIN B
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      0.7174 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5994 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      0.5826 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5148 LAYER met1 ;
    END A
    PIN GND
    END GND
END NOR2X1
MACRO NAND4BBXL
    PIN Y
        AntennaPartialMetalArea      1.4743 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1088 LAYER met1 ;
        AntennaDiffArea              1.1168 ;
    END Y
    PIN D
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.7555 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6966 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.6546 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5958 LAYER met1 ;
    END C
    PIN BN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8564 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7686 LAYER met1 ;
    END BN
    PIN AN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      1.0546 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8208 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NAND4BBXL
MACRO NAND4BBX4
    PIN Y
        AntennaPartialMetalArea      6.2950 LAYER met1 ;
        AntennaPartialMetalSideArea  4.4064 LAYER met1 ;
        AntennaDiffArea              5.3466 ;
    END Y
    PIN D
        AntennaGateArea              1.3752 ;
        AntennaPartialMetalArea      4.5876 LAYER met1 ;
        AntennaPartialMetalSideArea  3.5550 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              1.3752 ;
        AntennaPartialMetalArea      4.2958 LAYER met1 ;
        AntennaPartialMetalSideArea  3.5190 LAYER met1 ;
    END C
    PIN BN
        AntennaGateArea              0.5508 ;
        AntennaPartialMetalArea      0.7872 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5868 LAYER met1 ;
    END BN
    PIN AN
        AntennaGateArea              0.5508 ;
        AntennaPartialMetalArea      0.7807 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5976 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NAND4BBX4
MACRO NAND4BBX2
    PIN Y
        AntennaPartialMetalArea      3.0615 LAYER met1 ;
        AntennaPartialMetalSideArea  2.3310 LAYER met1 ;
        AntennaDiffArea              2.7144 ;
    END Y
    PIN D
        AntennaGateArea              0.7020 ;
        AntennaPartialMetalArea      2.4673 LAYER met1 ;
        AntennaPartialMetalSideArea  2.0736 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.7020 ;
        AntennaPartialMetalArea      1.9576 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6290 LAYER met1 ;
    END C
    PIN BN
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.7073 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6318 LAYER met1 ;
    END BN
    PIN AN
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.6780 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5904 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NAND4BBX2
MACRO NAND4BBX1
    PIN Y
        AntennaPartialMetalArea      1.4787 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1070 LAYER met1 ;
        AntennaDiffArea              1.5614 ;
    END Y
    PIN D
        AntennaGateArea              0.3456 ;
        AntennaPartialMetalArea      0.7417 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6696 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.3456 ;
        AntennaPartialMetalArea      0.6060 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5472 LAYER met1 ;
    END C
    PIN BN
        AntennaGateArea              0.1332 ;
        AntennaPartialMetalArea      0.8768 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8010 LAYER met1 ;
    END BN
    PIN AN
        AntennaGateArea              0.1332 ;
        AntennaPartialMetalArea      0.9840 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7902 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NAND4BBX1
MACRO NAND4BXL
    PIN Y
        AntennaPartialMetalArea      1.5783 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0926 LAYER met1 ;
        AntennaDiffArea              1.1000 ;
    END Y
    PIN D
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.6797 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5850 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.6226 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5706 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.7985 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6696 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7738 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6372 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NAND4BXL
MACRO NAND4BX4
    PIN Y
        AntennaPartialMetalArea      5.3460 LAYER met1 ;
        AntennaPartialMetalSideArea  3.7296 LAYER met1 ;
        AntennaDiffArea              5.3070 ;
    END Y
    PIN D
        AntennaGateArea              1.3752 ;
        AntennaPartialMetalArea      4.2823 LAYER met1 ;
        AntennaPartialMetalSideArea  3.4074 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              1.3752 ;
        AntennaPartialMetalArea      4.5573 LAYER met1 ;
        AntennaPartialMetalSideArea  3.5460 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              1.3752 ;
        AntennaPartialMetalArea      3.4770 LAYER met1 ;
        AntennaPartialMetalSideArea  2.8008 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.5508 ;
        AntennaPartialMetalArea      0.8207 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6120 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NAND4BX4
MACRO NAND4BX2
    PIN Y
        AntennaPartialMetalArea      2.4150 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8378 LAYER met1 ;
        AntennaDiffArea              2.7144 ;
    END Y
    PIN D
        AntennaGateArea              0.7020 ;
        AntennaPartialMetalArea      2.4673 LAYER met1 ;
        AntennaPartialMetalSideArea  2.0736 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.7020 ;
        AntennaPartialMetalArea      1.9841 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6398 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.7020 ;
        AntennaPartialMetalArea      1.4389 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2006 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.6780 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5904 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NAND4BX2
MACRO NAND4BX1
    PIN Y
        AntennaPartialMetalArea      1.5906 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0998 LAYER met1 ;
        AntennaDiffArea              1.4856 ;
    END Y
    PIN D
        AntennaGateArea              0.3456 ;
        AntennaPartialMetalArea      0.6582 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5814 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.3456 ;
        AntennaPartialMetalArea      0.6257 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5724 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.3456 ;
        AntennaPartialMetalArea      0.8246 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6768 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.1332 ;
        AntennaPartialMetalArea      0.7470 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6534 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NAND4BX1
MACRO NAND4XL
    PIN Y
        AntennaPartialMetalArea      1.5834 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1700 LAYER met1 ;
        AntennaDiffArea              1.1000 ;
    END Y
    PIN D
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.9031 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6732 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.6863 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6030 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.6550 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5886 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.7748 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6930 LAYER met1 ;
    END A
    PIN GND
    END GND
END NAND4XL
MACRO NAND4X4
    PIN Y
        AntennaPartialMetalArea      5.1796 LAYER met1 ;
        AntennaPartialMetalSideArea  3.6216 LAYER met1 ;
        AntennaDiffArea              5.3478 ;
    END Y
    PIN D
        AntennaGateArea              1.3752 ;
        AntennaPartialMetalArea      4.4517 LAYER met1 ;
        AntennaPartialMetalSideArea  3.3516 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              1.3752 ;
        AntennaPartialMetalArea      4.4144 LAYER met1 ;
        AntennaPartialMetalSideArea  3.5460 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              1.3752 ;
        AntennaPartialMetalArea      3.5375 LAYER met1 ;
        AntennaPartialMetalSideArea  2.8386 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              1.3752 ;
        AntennaPartialMetalArea      2.1485 LAYER met1 ;
        AntennaPartialMetalSideArea  2.0556 LAYER met1 ;
    END A
    PIN GND
    END GND
END NAND4X4
MACRO NAND4X2
    PIN Y
        AntennaPartialMetalArea      2.5632 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9260 LAYER met1 ;
        AntennaDiffArea              2.7144 ;
    END Y
    PIN D
        AntennaGateArea              0.7020 ;
        AntennaPartialMetalArea      2.4945 LAYER met1 ;
        AntennaPartialMetalSideArea  2.0160 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.7020 ;
        AntennaPartialMetalArea      1.9288 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6128 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.7020 ;
        AntennaPartialMetalArea      1.3986 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2060 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.7020 ;
        AntennaPartialMetalArea      0.9681 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8730 LAYER met1 ;
    END A
    PIN GND
    END GND
END NAND4X2
MACRO NAND4X1
    PIN Y
        AntennaPartialMetalArea      1.5815 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1700 LAYER met1 ;
        AntennaDiffArea              1.4856 ;
    END Y
    PIN D
        AntennaGateArea              0.3456 ;
        AntennaPartialMetalArea      0.9271 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6786 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.3456 ;
        AntennaPartialMetalArea      0.6863 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6030 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.3456 ;
        AntennaPartialMetalArea      0.6550 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5886 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.3456 ;
        AntennaPartialMetalArea      0.7773 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6894 LAYER met1 ;
    END A
    PIN GND
    END GND
END NAND4X1
MACRO NAND3BXL
    PIN Y
        AntennaPartialMetalArea      1.5723 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0440 LAYER met1 ;
        AntennaDiffArea              1.4184 ;
    END Y
    PIN C
        AntennaGateArea              0.2340 ;
        AntennaPartialMetalArea      1.0544 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0080 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.2340 ;
        AntennaPartialMetalArea      0.6902 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6264 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8072 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7470 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NAND3BXL
MACRO NAND3BX4
    PIN Y
        AntennaPartialMetalArea      5.5156 LAYER met1 ;
        AntennaPartialMetalSideArea  2.9916 LAYER met1 ;
        AntennaDiffArea              5.0720 ;
    END Y
    PIN C
        AntennaGateArea              1.2960 ;
        AntennaPartialMetalArea      2.6171 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2014 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              1.2960 ;
        AntennaPartialMetalArea      2.7293 LAYER met1 ;
        AntennaPartialMetalSideArea  2.3616 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.5040 ;
        AntennaPartialMetalArea      0.6931 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5922 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NAND3BX4
MACRO NAND3BX2
    PIN Y
        AntennaPartialMetalArea      1.9488 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4850 LAYER met1 ;
        AntennaDiffArea              2.5368 ;
    END Y
    PIN C
        AntennaGateArea              0.6696 ;
        AntennaPartialMetalArea      2.0313 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6452 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.6696 ;
        AntennaPartialMetalArea      1.4526 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2258 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.7226 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6444 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NAND3BX2
MACRO NAND3BX1
    PIN Y
        AntennaPartialMetalArea      1.2192 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9126 LAYER met1 ;
        AntennaDiffArea              1.5168 ;
    END Y
    PIN C
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7490 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6660 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7168 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6300 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.1332 ;
        AntennaPartialMetalArea      0.7175 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6408 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NAND3BX1
MACRO NAND3XL
    PIN Y
        AntennaPartialMetalArea      1.5849 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0548 LAYER met1 ;
        AntennaDiffArea              1.4120 ;
    END Y
    PIN C
        AntennaGateArea              0.2340 ;
        AntennaPartialMetalArea      1.2338 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1304 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.2340 ;
        AntennaPartialMetalArea      0.6942 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6336 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.2340 ;
        AntennaPartialMetalArea      0.6744 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6120 LAYER met1 ;
    END A
    PIN GND
    END GND
END NAND3XL
MACRO NAND3X4
    PIN Y
        AntennaPartialMetalArea      5.0487 LAYER met1 ;
        AntennaPartialMetalSideArea  3.0348 LAYER met1 ;
        AntennaDiffArea              5.0842 ;
    END Y
    PIN C
        AntennaGateArea              1.2960 ;
        AntennaPartialMetalArea      2.6298 LAYER met1 ;
        AntennaPartialMetalSideArea  2.1942 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              1.2960 ;
        AntennaPartialMetalArea      2.7308 LAYER met1 ;
        AntennaPartialMetalSideArea  2.3670 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              1.2960 ;
        AntennaPartialMetalArea      2.5232 LAYER met1 ;
        AntennaPartialMetalSideArea  2.1222 LAYER met1 ;
    END A
    PIN GND
    END GND
END NAND3X4
MACRO NAND3X2
    PIN Y
        AntennaPartialMetalArea      1.5614 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0656 LAYER met1 ;
        AntennaDiffArea              2.5924 ;
    END Y
    PIN C
        AntennaGateArea              0.6732 ;
        AntennaPartialMetalArea      2.5638 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9602 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.6732 ;
        AntennaPartialMetalArea      1.2967 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1160 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.6732 ;
        AntennaPartialMetalArea      0.7397 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6624 LAYER met1 ;
    END A
    PIN GND
    END GND
END NAND3X2
MACRO NAND3X1
    PIN Y
        AntennaPartialMetalArea      1.6308 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9720 LAYER met1 ;
        AntennaDiffArea              1.5384 ;
    END Y
    PIN C
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7617 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6858 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7231 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6444 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.8180 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7434 LAYER met1 ;
    END A
    PIN GND
    END GND
END NAND3X1
MACRO NAND2BXL
    PIN Y
        AntennaPartialMetalArea      1.0272 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7524 LAYER met1 ;
        AntennaDiffArea              0.6624 ;
    END Y
    PIN B
        AntennaGateArea              0.2160 ;
        AntennaPartialMetalArea      0.7157 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6408 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7172 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6282 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NAND2BXL
MACRO NAND2BX4
    PIN Y
        AntennaPartialMetalArea      3.0695 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8522 LAYER met1 ;
        AntennaDiffArea              3.2076 ;
    END Y
    PIN B
        AntennaGateArea              1.2276 ;
        AntennaPartialMetalArea      1.8245 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5354 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.4860 ;
        AntennaPartialMetalArea      0.8521 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6516 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NAND2BX4
MACRO NAND2BX2
    PIN Y
        AntennaPartialMetalArea      1.3450 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0512 LAYER met1 ;
        AntennaDiffArea              1.4622 ;
    END Y
    PIN B
        AntennaGateArea              0.6336 ;
        AntennaPartialMetalArea      1.5382 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3014 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.2412 ;
        AntennaPartialMetalArea      0.7748 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6480 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NAND2BX2
MACRO NAND2BX1
    PIN Y
        AntennaPartialMetalArea      1.1148 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7956 LAYER met1 ;
        AntennaDiffArea              0.9380 ;
    END Y
    PIN B
        AntennaGateArea              0.3060 ;
        AntennaPartialMetalArea      0.6635 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5886 LAYER met1 ;
    END B
    PIN AN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6139 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5490 LAYER met1 ;
    END AN
    PIN GND
    END GND
END NAND2BX1
MACRO NAND2XL
    PIN Y
        AntennaPartialMetalArea      0.9930 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6426 LAYER met1 ;
        AntennaDiffArea              0.6848 ;
    END Y
    PIN B
        AntennaGateArea              0.2160 ;
        AntennaPartialMetalArea      0.7301 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6300 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.2160 ;
        AntennaPartialMetalArea      0.7133 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6444 LAYER met1 ;
    END A
    PIN GND
    END GND
END NAND2XL
MACRO NAND2X4
    PIN Y
        AntennaPartialMetalArea      3.0803 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9188 LAYER met1 ;
        AntennaDiffArea              3.2160 ;
    END Y
    PIN B
        AntennaGateArea              1.2276 ;
        AntennaPartialMetalArea      2.2497 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5786 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              1.2276 ;
        AntennaPartialMetalArea      1.9082 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6002 LAYER met1 ;
    END A
    PIN GND
    END GND
END NAND2X4
MACRO NAND2X2
    PIN Y
        AntennaPartialMetalArea      1.5952 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1250 LAYER met1 ;
        AntennaDiffArea              1.4278 ;
    END Y
    PIN B
        AntennaGateArea              0.6336 ;
        AntennaPartialMetalArea      1.6049 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3356 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.6336 ;
        AntennaPartialMetalArea      1.0374 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9018 LAYER met1 ;
    END A
    PIN GND
    END GND
END NAND2X2
MACRO NAND2X1
    PIN Y
        AntennaPartialMetalArea      0.8886 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6192 LAYER met1 ;
        AntennaDiffArea              0.9198 ;
    END Y
    PIN B
        AntennaGateArea              0.3024 ;
        AntennaPartialMetalArea      0.6304 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5454 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.3024 ;
        AntennaPartialMetalArea      0.5920 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5166 LAYER met1 ;
    END A
    PIN GND
    END GND
END NAND2X1
MACRO MXI4XL
    PIN Y
        AntennaPartialMetalArea      1.0654 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7974 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END Y
    PIN S1
        AntennaGateArea              0.3816 ;
        AntennaPartialMetalArea      2.0676 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9890 LAYER met1 ;
    END S1
    PIN S0
        AntennaGateArea              0.6336 ;
        AntennaPartialMetalArea      3.3944 LAYER met1 ;
        AntennaPartialMetalSideArea  3.3012 LAYER met1 ;
    END S0
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7920 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6498 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7320 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6372 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6454 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5688 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8448 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6444 LAYER met1 ;
    END A
    PIN GND
    END GND
END MXI4XL
MACRO MXI4X4
    PIN Y
        AntennaPartialMetalArea      1.3526 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6894 LAYER met1 ;
        AntennaDiffArea              1.7400 ;
    END Y
    PIN S1
        AntennaGateArea              0.7380 ;
        AntennaPartialMetalArea      1.6766 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5912 LAYER met1 ;
    END S1
    PIN S0
        AntennaGateArea              1.2060 ;
        AntennaPartialMetalArea      3.0174 LAYER met1 ;
        AntennaPartialMetalSideArea  2.9538 LAYER met1 ;
    END S0
    PIN D
        AntennaGateArea              0.4284 ;
        AntennaPartialMetalArea      0.8073 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5832 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.4320 ;
        AntennaPartialMetalArea      0.7652 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6516 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.4284 ;
        AntennaPartialMetalArea      0.6660 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5940 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.4320 ;
        AntennaPartialMetalArea      0.8101 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5994 LAYER met1 ;
    END A
    PIN GND
    END GND
END MXI4X4
MACRO MXI4X2
    PIN Y
        AntennaPartialMetalArea      0.8597 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6174 LAYER met1 ;
        AntennaDiffArea              1.5768 ;
    END Y
    PIN S1
        AntennaGateArea              0.6012 ;
        AntennaPartialMetalArea      1.7756 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6596 LAYER met1 ;
    END S1
    PIN S0
        AntennaGateArea              0.9540 ;
        AntennaPartialMetalArea      3.1704 LAYER met1 ;
        AntennaPartialMetalSideArea  3.0870 LAYER met1 ;
    END S0
    PIN D
        AntennaGateArea              0.3312 ;
        AntennaPartialMetalArea      0.7819 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6318 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.3420 ;
        AntennaPartialMetalArea      0.8084 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6948 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.3420 ;
        AntennaPartialMetalArea      0.6660 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6048 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.3420 ;
        AntennaPartialMetalArea      0.8525 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6336 LAYER met1 ;
    END A
    PIN GND
    END GND
END MXI4X2
MACRO MXI4X1
    PIN Y
        AntennaPartialMetalArea      0.9122 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5544 LAYER met1 ;
        AntennaDiffArea              0.7740 ;
    END Y
    PIN S1
        AntennaGateArea              0.3456 ;
        AntennaPartialMetalArea      2.1182 LAYER met1 ;
        AntennaPartialMetalSideArea  2.0340 LAYER met1 ;
    END S1
    PIN S0
        AntennaGateArea              0.4716 ;
        AntennaPartialMetalArea      3.5979 LAYER met1 ;
        AntennaPartialMetalSideArea  3.4974 LAYER met1 ;
    END S0
    PIN D
        AntennaGateArea              0.1692 ;
        AntennaPartialMetalArea      0.7428 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6012 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.1692 ;
        AntennaPartialMetalArea      0.6722 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6246 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.1692 ;
        AntennaPartialMetalArea      0.7374 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6408 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.1692 ;
        AntennaPartialMetalArea      0.9882 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8010 LAYER met1 ;
    END A
    PIN GND
    END GND
END MXI4X1
MACRO MXI2XL
    PIN Y
        AntennaPartialMetalArea      0.6782 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4698 LAYER met1 ;
        AntennaDiffArea              0.8456 ;
    END Y
    PIN S0
        AntennaGateArea              0.3816 ;
        AntennaPartialMetalArea      2.0528 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9818 LAYER met1 ;
    END S0
    PIN B
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6668 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5850 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.6614 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5634 LAYER met1 ;
    END A
    PIN GND
    END GND
END MXI2XL
MACRO MXI2X4
    PIN Y
        AntennaPartialMetalArea      3.0987 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8414 LAYER met1 ;
        AntennaDiffArea              4.9690 ;
    END Y
    PIN S0
        AntennaGateArea              1.5552 ;
        AntennaPartialMetalArea      3.5302 LAYER met1 ;
        AntennaPartialMetalSideArea  2.8836 LAYER met1 ;
    END S0
    PIN B
        AntennaGateArea              1.1088 ;
        AntennaPartialMetalArea      1.0914 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8028 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              1.1088 ;
        AntennaPartialMetalArea      1.2424 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8838 LAYER met1 ;
    END A
    PIN GND
    END GND
END MXI2X4
MACRO MXI2X2
    PIN Y
        AntennaPartialMetalArea      0.7892 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6120 LAYER met1 ;
        AntennaDiffArea              1.8596 ;
    END Y
    PIN S0
        AntennaGateArea              0.7308 ;
        AntennaPartialMetalArea      1.6674 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5894 LAYER met1 ;
    END S0
    PIN B
        AntennaGateArea              0.5076 ;
        AntennaPartialMetalArea      0.6740 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5706 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5496 ;
        AntennaPartialMetalArea      0.7256 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6048 LAYER met1 ;
    END A
    PIN GND
    END GND
END MXI2X2
MACRO MXI2X1
    PIN Y
        AntennaPartialMetalArea      0.6782 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4698 LAYER met1 ;
        AntennaDiffArea              1.0028 ;
    END Y
    PIN S0
        AntennaGateArea              0.4356 ;
        AntennaPartialMetalArea      2.0822 LAYER met1 ;
        AntennaPartialMetalSideArea  2.0034 LAYER met1 ;
    END S0
    PIN B
        AntennaGateArea              0.2988 ;
        AntennaPartialMetalArea      0.6164 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5346 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.2988 ;
        AntennaPartialMetalArea      0.6540 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5544 LAYER met1 ;
    END A
    PIN GND
    END GND
END MXI2X1
MACRO MX4XL
    PIN Y
        AntennaPartialMetalArea      1.0202 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6030 LAYER met1 ;
        AntennaDiffArea              0.6609 ;
    END Y
    PIN S1
        AntennaGateArea              0.3816 ;
        AntennaPartialMetalArea      1.7000 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5858 LAYER met1 ;
    END S1
    PIN S0
        AntennaGateArea              0.6336 ;
        AntennaPartialMetalArea      3.4052 LAYER met1 ;
        AntennaPartialMetalSideArea  3.3120 LAYER met1 ;
    END S0
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6454 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5688 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8424 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6498 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7920 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6498 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7639 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6156 LAYER met1 ;
    END A
    PIN GND
    END GND
END MX4XL
MACRO MX4X4
    PIN Y
        AntennaPartialMetalArea      1.0934 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5418 LAYER met1 ;
        AntennaDiffArea              1.4682 ;
    END Y
    PIN S1
        AntennaGateArea              0.7560 ;
        AntennaPartialMetalArea      2.6261 LAYER met1 ;
        AntennaPartialMetalSideArea  2.1312 LAYER met1 ;
    END S1
    PIN S0
        AntennaGateArea              1.4868 ;
        AntennaPartialMetalArea      5.3448 LAYER met1 ;
        AntennaPartialMetalSideArea  4.5072 LAYER met1 ;
    END S0
    PIN D
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.6184 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5652 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.7519 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5778 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.5882 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5184 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.5924 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5238 LAYER met1 ;
    END A
    PIN GND
    END GND
END MX4X4
MACRO MX4X2
    PIN Y
        AntennaPartialMetalArea      1.0364 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6804 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Y
    PIN S1
        AntennaGateArea              0.7560 ;
        AntennaPartialMetalArea      2.6151 LAYER met1 ;
        AntennaPartialMetalSideArea  2.1186 LAYER met1 ;
    END S1
    PIN S0
        AntennaGateArea              1.4868 ;
        AntennaPartialMetalArea      5.4419 LAYER met1 ;
        AntennaPartialMetalSideArea  4.6044 LAYER met1 ;
    END S0
    PIN D
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.6184 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5652 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.7230 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5814 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.5882 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5184 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.5924 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5238 LAYER met1 ;
    END A
    PIN GND
    END GND
END MX4X2
MACRO MX4X1
    PIN Y
        AntennaPartialMetalArea      1.0250 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7002 LAYER met1 ;
        AntennaDiffArea              0.7768 ;
    END Y
    PIN S1
        AntennaGateArea              0.4536 ;
        AntennaPartialMetalArea      1.6446 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5804 LAYER met1 ;
    END S1
    PIN S0
        AntennaGateArea              0.9108 ;
        AntennaPartialMetalArea      3.2432 LAYER met1 ;
        AntennaPartialMetalSideArea  3.1500 LAYER met1 ;
    END S0
    PIN D
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      0.6250 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5634 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      0.7525 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6192 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      0.7789 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6210 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      0.7346 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5850 LAYER met1 ;
    END A
    PIN GND
    END GND
END MX4X1
MACRO MX2XL
    PIN Y
        AntennaPartialMetalArea      0.8834 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6516 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END Y
    PIN S0
        AntennaGateArea              0.3816 ;
        AntennaPartialMetalArea      1.9570 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8846 LAYER met1 ;
    END S0
    PIN B
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8267 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7200 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6876 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6120 LAYER met1 ;
    END A
    PIN GND
    END GND
END MX2XL
MACRO MX2X4
    PIN Y
        AntennaPartialMetalArea      1.5300 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9774 LAYER met1 ;
        AntennaDiffArea              1.5629 ;
    END Y
    PIN S0
        AntennaGateArea              0.7488 ;
        AntennaPartialMetalArea      1.7108 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6416 LAYER met1 ;
    END S0
    PIN B
        AntennaGateArea              0.4932 ;
        AntennaPartialMetalArea      0.6376 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5256 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5472 ;
        AntennaPartialMetalArea      0.6360 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5652 LAYER met1 ;
    END A
    PIN GND
    END GND
END MX2X4
MACRO MX2X2
    PIN Y
        AntennaPartialMetalArea      1.0416 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6912 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Y
    PIN S0
        AntennaGateArea              0.6012 ;
        AntennaPartialMetalArea      2.1421 LAYER met1 ;
        AntennaPartialMetalSideArea  2.0286 LAYER met1 ;
    END S0
    PIN B
        AntennaGateArea              0.4248 ;
        AntennaPartialMetalArea      0.7248 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5886 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.4320 ;
        AntennaPartialMetalArea      0.7138 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6354 LAYER met1 ;
    END A
    PIN GND
    END GND
END MX2X2
MACRO MX2X1
    PIN Y
        AntennaPartialMetalArea      0.8514 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6318 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Y
    PIN S0
        AntennaGateArea              0.3456 ;
        AntennaPartialMetalArea      1.9248 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8522 LAYER met1 ;
    END S0
    PIN B
        AntennaGateArea              0.2160 ;
        AntennaPartialMetalArea      0.8319 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7254 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.2160 ;
        AntennaPartialMetalArea      0.7196 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6318 LAYER met1 ;
    END A
    PIN GND
    END GND
END MX2X1
MACRO JKFFSRXL
    PIN SN
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      2.1914 LAYER met1 ;
        AntennaPartialMetalSideArea  2.1186 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      1.0489 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8640 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.3861 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0584 LAYER met1 ;
        AntennaDiffArea              0.6081 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6508 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4644 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END Q
    PIN K
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.8073 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7650 LAYER met1 ;
    END K
    PIN J
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.7977 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6714 LAYER met1 ;
    END J
    PIN CK
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6104 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5436 LAYER met1 ;
    END CK
    PIN GND
    END GND
END JKFFSRXL
MACRO JKFFSRX4
    PIN SN
        AntennaGateArea              0.5688 ;
        AntennaPartialMetalArea      1.8384 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7712 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      1.1532 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9000 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.3094 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6318 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.5202 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6714 LAYER met1 ;
        AntennaDiffArea              1.4562 ;
    END Q
    PIN K
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.8140 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7740 LAYER met1 ;
    END K
    PIN J
        AntennaGateArea              0.1260 ;
        AntennaPartialMetalArea      0.6895 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6390 LAYER met1 ;
    END J
    PIN CK
        AntennaGateArea              0.2052 ;
        AntennaPartialMetalArea      0.5979 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5346 LAYER met1 ;
    END CK
    PIN GND
    END GND
END JKFFSRX4
MACRO JKFFSRX2
    PIN SN
        AntennaGateArea              0.5688 ;
        AntennaPartialMetalArea      1.8384 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7712 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      1.1532 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9000 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.7612 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5724 LAYER met1 ;
        AntennaDiffArea              1.3938 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.0830 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7272 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Q
    PIN K
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.8140 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7740 LAYER met1 ;
    END K
    PIN J
        AntennaGateArea              0.1260 ;
        AntennaPartialMetalArea      0.6895 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6390 LAYER met1 ;
    END J
    PIN CK
        AntennaGateArea              0.2052 ;
        AntennaPartialMetalArea      0.5979 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5346 LAYER met1 ;
    END CK
    PIN GND
    END GND
END JKFFSRX2
MACRO JKFFSRX1
    PIN SN
        AntennaGateArea              0.3492 ;
        AntennaPartialMetalArea      2.1444 LAYER met1 ;
        AntennaPartialMetalSideArea  2.0772 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.1620 ;
        AntennaPartialMetalArea      1.0372 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8532 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.4293 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0908 LAYER met1 ;
        AntennaDiffArea              0.8101 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6410 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4572 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN K
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.8140 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7740 LAYER met1 ;
    END K
    PIN J
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      0.6895 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6390 LAYER met1 ;
    END J
    PIN CK
        AntennaGateArea              0.1692 ;
        AntennaPartialMetalArea      0.5979 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5346 LAYER met1 ;
    END CK
    PIN GND
    END GND
END JKFFSRX1
MACRO JKFFSXL
    PIN SN
        AntennaGateArea              0.2808 ;
        AntennaPartialMetalArea      3.0315 LAYER met1 ;
        AntennaPartialMetalSideArea  2.4966 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      0.7396 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5436 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6332 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4590 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END Q
    PIN K
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.6687 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5940 LAYER met1 ;
    END K
    PIN J
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.6869 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6174 LAYER met1 ;
    END J
    PIN CK
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.6082 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5436 LAYER met1 ;
    END CK
    PIN GND
    END GND
END JKFFSXL
MACRO JKFFSX4
    PIN SN
        AntennaGateArea              0.9648 ;
        AntennaPartialMetalArea      4.6147 LAYER met1 ;
        AntennaPartialMetalSideArea  3.7818 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      1.0686 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4644 LAYER met1 ;
        AntennaDiffArea              1.4562 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.1665 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5022 LAYER met1 ;
        AntennaDiffArea              1.4562 ;
    END Q
    PIN K
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.6868 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6084 LAYER met1 ;
    END K
    PIN J
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7291 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6642 LAYER met1 ;
    END J
    PIN CK
        AntennaGateArea              0.2628 ;
        AntennaPartialMetalArea      0.5830 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5058 LAYER met1 ;
    END CK
    PIN GND
    END GND
END JKFFSX4
MACRO JKFFSX2
    PIN SN
        AntennaGateArea              0.5436 ;
        AntennaPartialMetalArea      3.3996 LAYER met1 ;
        AntennaPartialMetalSideArea  2.8188 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      0.7179 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4860 LAYER met1 ;
        AntennaDiffArea              1.1455 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.7704 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5670 LAYER met1 ;
        AntennaDiffArea              1.1879 ;
    END Q
    PIN K
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.6687 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5940 LAYER met1 ;
    END K
    PIN J
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      0.7229 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6534 LAYER met1 ;
    END J
    PIN CK
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.6082 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5436 LAYER met1 ;
    END CK
    PIN GND
    END GND
END JKFFSX2
MACRO JKFFSX1
    PIN SN
        AntennaGateArea              0.3744 ;
        AntennaPartialMetalArea      2.9577 LAYER met1 ;
        AntennaPartialMetalSideArea  2.4228 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      0.7332 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5400 LAYER met1 ;
        AntennaDiffArea              0.7488 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6588 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4698 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN K
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.6687 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5940 LAYER met1 ;
    END K
    PIN J
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      0.7229 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6534 LAYER met1 ;
    END J
    PIN CK
        AntennaGateArea              0.1692 ;
        AntennaPartialMetalArea      0.6082 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5436 LAYER met1 ;
    END CK
    PIN GND
    END GND
END JKFFSX1
MACRO JKFFRXL
    PIN RN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7850 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7218 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.8800 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6786 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.7412 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5490 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END Q
    PIN K
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.6352 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5958 LAYER met1 ;
    END K
    PIN J
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.7298 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6516 LAYER met1 ;
    END J
    PIN CK
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.6556 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5670 LAYER met1 ;
    END CK
    PIN GND
    END GND
END JKFFRXL
MACRO JKFFRX4
    PIN RN
        AntennaGateArea              0.4176 ;
        AntennaPartialMetalArea      0.9312 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7272 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.9611 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4860 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.9160 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4662 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END Q
    PIN K
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.6768 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6174 LAYER met1 ;
    END K
    PIN J
        AntennaGateArea              0.1620 ;
        AntennaPartialMetalArea      0.7498 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6768 LAYER met1 ;
    END J
    PIN CK
        AntennaGateArea              0.2988 ;
        AntennaPartialMetalArea      0.6160 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5274 LAYER met1 ;
    END CK
    PIN GND
    END GND
END JKFFRX4
MACRO JKFFRX2
    PIN RN
        AntennaGateArea              0.2340 ;
        AntennaPartialMetalArea      0.5807 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5202 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.6968 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4824 LAYER met1 ;
        AntennaDiffArea              1.1879 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8278 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6012 LAYER met1 ;
        AntennaDiffArea              1.1879 ;
    END Q
    PIN K
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.6374 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5958 LAYER met1 ;
    END K
    PIN J
        AntennaGateArea              0.1116 ;
        AntennaPartialMetalArea      0.7642 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6912 LAYER met1 ;
    END J
    PIN CK
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.6394 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5508 LAYER met1 ;
    END CK
    PIN GND
    END GND
END JKFFRX2
MACRO JKFFRX1
    PIN RN
        AntennaGateArea              0.1620 ;
        AntennaPartialMetalArea      0.7616 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6984 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.8695 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6696 LAYER met1 ;
        AntennaDiffArea              0.7200 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.7436 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5508 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN K
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.6542 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6102 LAYER met1 ;
    END K
    PIN J
        AntennaGateArea              0.1116 ;
        AntennaPartialMetalArea      0.7642 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6912 LAYER met1 ;
    END J
    PIN CK
        AntennaGateArea              0.1692 ;
        AntennaPartialMetalArea      0.6466 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5580 LAYER met1 ;
    END CK
    PIN GND
    END GND
END JKFFRX1
MACRO JKFFXL
    PIN QN
        AntennaPartialMetalArea      0.6192 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4662 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6286 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4320 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END Q
    PIN K
        AntennaGateArea              0.2016 ;
        AntennaPartialMetalArea      0.6777 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6354 LAYER met1 ;
    END K
    PIN J
        AntennaGateArea              0.1404 ;
        AntennaPartialMetalArea      0.7491 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6606 LAYER met1 ;
    END J
    PIN CK
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8250 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6876 LAYER met1 ;
    END CK
    PIN GND
    END GND
END JKFFXL
MACRO JKFFX4
    PIN QN
        AntennaPartialMetalArea      0.9409 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4392 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.9800 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4770 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END Q
    PIN K
        AntennaGateArea              0.2592 ;
        AntennaPartialMetalArea      0.6207 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5832 LAYER met1 ;
    END K
    PIN J
        AntennaGateArea              0.1116 ;
        AntennaPartialMetalArea      0.7935 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7200 LAYER met1 ;
    END J
    PIN CK
        AntennaGateArea              0.5544 ;
        AntennaPartialMetalArea      0.6080 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5310 LAYER met1 ;
    END CK
    PIN GND
    END GND
END JKFFX4
MACRO JKFFX2
    PIN QN
        AntennaPartialMetalArea      0.7487 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5454 LAYER met1 ;
        AntennaDiffArea              1.4215 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8372 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6192 LAYER met1 ;
        AntennaDiffArea              1.4095 ;
    END Q
    PIN K
        AntennaGateArea              0.1404 ;
        AntennaPartialMetalArea      0.7280 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6732 LAYER met1 ;
    END K
    PIN J
        AntennaGateArea              0.1116 ;
        AntennaPartialMetalArea      1.0380 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9486 LAYER met1 ;
    END J
    PIN CK
        AntennaGateArea              0.3024 ;
        AntennaPartialMetalArea      0.7503 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6606 LAYER met1 ;
    END CK
    PIN GND
    END GND
END JKFFX2
MACRO JKFFX1
    PIN QN
        AntennaPartialMetalArea      1.3708 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0314 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.7660 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4086 LAYER met1 ;
        AntennaDiffArea              0.7639 ;
    END Q
    PIN K
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      0.7373 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6786 LAYER met1 ;
    END K
    PIN J
        AntennaGateArea              0.1116 ;
        AntennaPartialMetalArea      0.7725 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6840 LAYER met1 ;
    END J
    PIN CK
        AntennaGateArea              0.2052 ;
        AntennaPartialMetalArea      0.7416 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6552 LAYER met1 ;
    END CK
    PIN GND
    END GND
END JKFFX1
MACRO INVXL
    PIN Y
        AntennaPartialMetalArea      0.5858 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4518 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END Y
    PIN A
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      1.0118 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8046 LAYER met1 ;
    END A
    PIN GND
    END GND
END INVXL
MACRO INVX8
    PIN Y
        AntennaPartialMetalArea      4.1472 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9486 LAYER met1 ;
        AntennaDiffArea              2.8704 ;
    END Y
    PIN A
        AntennaGateArea              2.2200 ;
        AntennaPartialMetalArea      2.3922 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6254 LAYER met1 ;
    END A
    PIN GND
    END GND
END INVX8
MACRO INVX4
    PIN Y
        AntennaPartialMetalArea      0.9228 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4806 LAYER met1 ;
        AntennaDiffArea              1.5345 ;
    END Y
    PIN A
        AntennaGateArea              1.0764 ;
        AntennaPartialMetalArea      1.3391 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9342 LAYER met1 ;
    END A
    PIN GND
    END GND
END INVX4
MACRO INVX3
    PIN Y
        AntennaPartialMetalArea      1.0983 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6192 LAYER met1 ;
        AntennaDiffArea              1.3224 ;
    END Y
    PIN A
        AntennaGateArea              0.8100 ;
        AntennaPartialMetalArea      1.1648 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8496 LAYER met1 ;
    END A
    PIN GND
    END GND
END INVX3
MACRO INVX2
    PIN Y
        AntennaPartialMetalArea      0.9431 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6282 LAYER met1 ;
        AntennaDiffArea              1.1100 ;
    END Y
    PIN A
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      1.3487 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9864 LAYER met1 ;
    END A
    PIN GND
    END GND
END INVX2
MACRO INVX20
    PIN Y
        AntennaPartialMetalArea      11.5662 LAYER met1 ;
        AntennaPartialMetalSideArea  2.6352 LAYER met1 ;
        AntennaDiffArea              7.8790 ;
    END Y
    PIN A
        AntennaGateArea              0.8682 ;
        AntennaPartialMetalArea      1.2720 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9000 LAYER met1 ;
    END A
    PIN GND
    END GND
END INVX20
MACRO INVX1
    PIN Y
        AntennaPartialMetalArea      0.6452 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4860 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Y
    PIN A
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.6740 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5760 LAYER met1 ;
    END A
    PIN GND
    END GND
END INVX1
MACRO INVX16
    PIN Y
        AntennaPartialMetalArea      10.3681 LAYER met1 ;
        AntennaPartialMetalSideArea  2.0880 LAYER met1 ;
        AntennaDiffArea              6.8783 ;
    END Y
    PIN A
        AntennaGateArea              0.6756 ;
        AntennaPartialMetalArea      0.9259 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7254 LAYER met1 ;
    END A
    PIN GND
    END GND
END INVX16
MACRO INVX12
    PIN Y
        AntennaPartialMetalArea      6.8006 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4850 LAYER met1 ;
        AntennaDiffArea              4.5954 ;
    END Y
    PIN A
        AntennaGateArea              0.5298 ;
        AntennaPartialMetalArea      0.5768 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5166 LAYER met1 ;
    END A
    PIN GND
    END GND
END INVX12
MACRO HOLDX1
    PIN Y
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      1.7331 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4274 LAYER met1 ;
        AntennaDiffArea              0.4682 ;
    END Y
    PIN GND
    END GND
END HOLDX1
MACRO FILL8
    CLASS CORE SPACER ;
    PIN GND
    END GND
END FILL8
MACRO FILL64
    CLASS CORE SPACER ;
    PIN GND
    END GND
END FILL64
MACRO FILL4
    CLASS CORE SPACER ;
    PIN GND
    END GND
END FILL4
MACRO FILL32
    CLASS CORE SPACER ;
    PIN GND
    END GND
END FILL32
MACRO FILL2
    CLASS CORE SPACER ;
    PIN GND
    END GND
END FILL2
MACRO FILL16
    CLASS CORE SPACER ;
    PIN GND
    END GND
END FILL16
MACRO FILL1
    CLASS CORE SPACER ;
    PIN GND
    END GND
END FILL1
MACRO EDFFTRXL
    PIN RN
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      1.1926 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0548 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.7852 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6318 LAYER met1 ;
        AntennaDiffArea              0.6297 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.4770 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0620 LAYER met1 ;
        AntennaDiffArea              0.5628 ;
    END Q
    PIN E
        AntennaGateArea              0.3420 ;
        AntennaPartialMetalArea      2.2104 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7838 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.2052 ;
        AntennaPartialMetalArea      0.8779 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8082 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8493 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7326 LAYER met1 ;
    END CK
    PIN GND
    END GND
END EDFFTRXL
MACRO EDFFTRX4
    PIN RN
        AntennaGateArea              0.2412 ;
        AntennaPartialMetalArea      1.2141 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1160 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.0858 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5364 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.9595 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4788 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END Q
    PIN E
        AntennaGateArea              0.3924 ;
        AntennaPartialMetalArea      2.2659 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8450 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.2628 ;
        AntennaPartialMetalArea      0.9709 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9090 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.5436 ;
        AntennaPartialMetalArea      0.5672 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5148 LAYER met1 ;
    END CK
    PIN GND
    END GND
END EDFFTRX4
MACRO EDFFTRX2
    PIN RN
        AntennaGateArea              0.1332 ;
        AntennaPartialMetalArea      1.0638 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0026 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.0667 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8064 LAYER met1 ;
        AntennaDiffArea              1.3516 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.5536 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0962 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Q
    PIN E
        AntennaGateArea              0.2736 ;
        AntennaPartialMetalArea      2.1463 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8558 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.1440 ;
        AntennaPartialMetalArea      0.9882 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9036 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.3060 ;
        AntennaPartialMetalArea      0.8645 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7434 LAYER met1 ;
    END CK
    PIN GND
    END GND
END EDFFTRX2
MACRO EDFFTRX1
    PIN RN
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      1.0743 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0170 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.9085 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6642 LAYER met1 ;
        AntennaDiffArea              0.8668 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.3184 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9900 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN E
        AntennaGateArea              0.2376 ;
        AntennaPartialMetalArea      2.1195 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8396 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      0.9379 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8442 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2052 ;
        AntennaPartialMetalArea      0.8573 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7434 LAYER met1 ;
    END CK
    PIN GND
    END GND
END EDFFTRX1
MACRO EDFFXL
    PIN QN
        AntennaPartialMetalArea      0.6426 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4320 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.3668 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0332 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END Q
    PIN E
        AntennaGateArea              0.3276 ;
        AntennaPartialMetalArea      1.8462 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7280 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.7972 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7254 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.6511 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6120 LAYER met1 ;
    END CK
    PIN GND
    END GND
END EDFFXL
MACRO EDFFX4
    PIN QN
        AntennaPartialMetalArea      0.8877 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4536 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.9835 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4968 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END Q
    PIN E
        AntennaGateArea              0.3852 ;
        AntennaPartialMetalArea      1.8888 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7802 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.7438 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6642 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.5220 ;
        AntennaPartialMetalArea      0.6264 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5526 LAYER met1 ;
    END CK
    PIN GND
    END GND
END EDFFX4
MACRO EDFFX2
    PIN QN
        AntennaPartialMetalArea      0.7774 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5490 LAYER met1 ;
        AntennaDiffArea              1.2382 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.5064 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4212 LAYER met1 ;
        AntennaDiffArea              1.0530 ;
    END Q
    PIN E
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      1.7384 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6758 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.1404 ;
        AntennaPartialMetalArea      1.0423 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9342 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.3060 ;
        AntennaPartialMetalArea      0.6151 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5760 LAYER met1 ;
    END CK
    PIN GND
    END GND
END EDFFX2
MACRO EDFFX1
    PIN QN
        AntennaPartialMetalArea      0.6540 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4752 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.4020 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0548 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN E
        AntennaGateArea              0.2376 ;
        AntennaPartialMetalArea      1.8912 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7730 LAYER met1 ;
    END E
    PIN D
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      1.0332 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9072 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2052 ;
        AntennaPartialMetalArea      0.6271 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5850 LAYER met1 ;
    END CK
    PIN GND
    END GND
END EDFFX1
MACRO DLY4X1
    PIN Y
        AntennaPartialMetalArea      0.6572 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4734 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Y
    PIN A
        AntennaGateArea              0.1260 ;
        AntennaPartialMetalArea      0.6175 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5454 LAYER met1 ;
    END A
    PIN GND
    END GND
END DLY4X1
MACRO DLY3X1
    PIN Y
        AntennaPartialMetalArea      0.6572 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4734 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Y
    PIN A
        AntennaGateArea              0.1260 ;
        AntennaPartialMetalArea      0.6175 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5454 LAYER met1 ;
    END A
    PIN GND
    END GND
END DLY3X1
MACRO DLY2X1
    PIN Y
        AntennaPartialMetalArea      0.6572 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4734 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Y
    PIN A
        AntennaGateArea              0.1260 ;
        AntennaPartialMetalArea      0.6175 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5454 LAYER met1 ;
    END A
    PIN GND
    END GND
END DLY2X1
MACRO DLY1X1
    PIN Y
        AntennaPartialMetalArea      0.6572 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4734 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Y
    PIN A
        AntennaGateArea              0.1260 ;
        AntennaPartialMetalArea      0.6175 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5454 LAYER met1 ;
    END A
    PIN GND
    END GND
END DLY1X1
MACRO DFFTRXL
    PIN RN
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.6606 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5940 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.4786 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4014 LAYER met1 ;
        AntennaDiffArea              0.6250 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.3055 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9666 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END Q
    PIN D
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.7951 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7164 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6486 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5796 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFTRXL
MACRO DFFTRX4
    PIN RN
        AntennaGateArea              0.2124 ;
        AntennaPartialMetalArea      0.6739 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5814 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.8120 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4194 LAYER met1 ;
        AntennaDiffArea              1.4232 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.9478 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4716 LAYER met1 ;
        AntennaDiffArea              1.4232 ;
    END Q
    PIN D
        AntennaGateArea              0.2124 ;
        AntennaPartialMetalArea      0.8846 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8190 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.4932 ;
        AntennaPartialMetalArea      0.5610 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5094 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFTRX4
MACRO DFFTRX2
    PIN RN
        AntennaGateArea              0.1188 ;
        AntennaPartialMetalArea      0.6447 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5850 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.1338 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7596 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6826 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5310 LAYER met1 ;
        AntennaDiffArea              1.2292 ;
    END Q
    PIN D
        AntennaGateArea              0.1188 ;
        AntennaPartialMetalArea      0.7985 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7146 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      0.5684 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5076 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFTRX2
MACRO DFFTRX1
    PIN RN
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      0.6948 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6282 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.5564 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4554 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.3413 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9828 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN D
        AntennaGateArea              0.1080 ;
        AntennaPartialMetalArea      0.8095 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7308 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.6433 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6030 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFTRX1
MACRO DFFSRHQXL
    PIN SN
        AntennaGateArea              0.4968 ;
        AntennaPartialMetalArea      5.9024 LAYER met1 ;
        AntennaPartialMetalSideArea  4.6260 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6766 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6192 LAYER met1 ;
    END RN
    PIN Q
        AntennaPartialMetalArea      1.1558 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8712 LAYER met1 ;
        AntennaDiffArea              0.7760 ;
    END Q
    PIN D
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7710 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7074 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8173 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7488 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFSRHQXL
MACRO DFFSRHQX4
    PIN SN
        AntennaGateArea              1.7562 ;
        AntennaPartialMetalArea      7.3000 LAYER met1 ;
        AntennaPartialMetalSideArea  5.6736 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.8136 ;
        AntennaPartialMetalArea      1.3250 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9828 LAYER met1 ;
    END RN
    PIN Q
        AntennaPartialMetalArea      3.6826 LAYER met1 ;
        AntennaPartialMetalSideArea  2.3418 LAYER met1 ;
        AntennaDiffArea              4.8825 ;
    END Q
    PIN D
        AntennaGateArea              0.3960 ;
        AntennaPartialMetalArea      0.7027 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6264 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.5292 ;
        AntennaPartialMetalArea      0.6592 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5544 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFSRHQX4
MACRO DFFSRHQX2
    PIN SN
        AntennaGateArea              0.9720 ;
        AntennaPartialMetalArea      6.6418 LAYER met1 ;
        AntennaPartialMetalSideArea  5.0184 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.4428 ;
        AntennaPartialMetalArea      0.6858 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5796 LAYER met1 ;
    END RN
    PIN Q
        AntennaPartialMetalArea      1.8823 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2942 LAYER met1 ;
        AntennaDiffArea              2.5965 ;
    END Q
    PIN D
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      0.7410 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6930 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.3132 ;
        AntennaPartialMetalArea      0.6522 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5508 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFSRHQX2
MACRO DFFSRHQX1
    PIN SN
        AntennaGateArea              0.5688 ;
        AntennaPartialMetalArea      5.7096 LAYER met1 ;
        AntennaPartialMetalSideArea  4.5036 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7116 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6462 LAYER met1 ;
    END RN
    PIN Q
        AntennaPartialMetalArea      1.1464 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8802 LAYER met1 ;
        AntennaDiffArea              1.1060 ;
    END Q
    PIN D
        AntennaGateArea              0.1440 ;
        AntennaPartialMetalArea      0.7134 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5832 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2160 ;
        AntennaPartialMetalArea      0.6256 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5580 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFSRHQX1
MACRO DFFSRXL
    PIN SN
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      3.3297 LAYER met1 ;
        AntennaPartialMetalSideArea  2.7828 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7600 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6858 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.2484 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9324 LAYER met1 ;
        AntennaDiffArea              0.5849 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.4725 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7758 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END Q
    PIN D
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.7680 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6588 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.7606 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6858 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFSRXL
MACRO DFFSRX4
    PIN SN
        AntennaGateArea              0.9792 ;
        AntennaPartialMetalArea      4.4086 LAYER met1 ;
        AntennaPartialMetalSideArea  3.6414 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.4644 ;
        AntennaPartialMetalArea      0.6016 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5076 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.9768 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4338 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.2694 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4734 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END Q
    PIN D
        AntennaGateArea              0.2412 ;
        AntennaPartialMetalArea      0.7537 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6480 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.3132 ;
        AntennaPartialMetalArea      0.6239 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5706 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFSRX4
MACRO DFFSRX2
    PIN SN
        AntennaGateArea              0.5328 ;
        AntennaPartialMetalArea      3.1108 LAYER met1 ;
        AntennaPartialMetalSideArea  2.5362 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.8003 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7218 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.6387 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4734 LAYER met1 ;
        AntennaDiffArea              1.1363 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8068 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5922 LAYER met1 ;
        AntennaDiffArea              1.2341 ;
    END Q
    PIN D
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.6981 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6030 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.8243 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6552 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFSRX2
MACRO DFFSRX1
    PIN SN
        AntennaGateArea              0.3312 ;
        AntennaPartialMetalArea      3.2173 LAYER met1 ;
        AntennaPartialMetalSideArea  2.6514 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.8313 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7326 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.1636 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8964 LAYER met1 ;
        AntennaDiffArea              0.7743 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8177 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5976 LAYER met1 ;
        AntennaDiffArea              0.7740 ;
    END Q
    PIN D
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.6886 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5994 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.7181 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6174 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFSRX1
MACRO DFFSHQXL
    PIN SN
        AntennaGateArea              0.5112 ;
        AntennaPartialMetalArea      4.3824 LAYER met1 ;
        AntennaPartialMetalSideArea  3.3912 LAYER met1 ;
    END SN
    PIN Q
        AntennaPartialMetalArea      0.9094 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6912 LAYER met1 ;
        AntennaDiffArea              0.6624 ;
    END Q
    PIN D
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.9772 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8010 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.8777 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7488 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFSHQXL
MACRO DFFSHQX4
    PIN SN
        AntennaGateArea              1.7028 ;
        AntennaPartialMetalArea      6.4089 LAYER met1 ;
        AntennaPartialMetalSideArea  4.6026 LAYER met1 ;
    END SN
    PIN Q
        AntennaPartialMetalArea      3.0963 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8090 LAYER met1 ;
        AntennaDiffArea              3.2540 ;
    END Q
    PIN D
        AntennaGateArea              0.2988 ;
        AntennaPartialMetalArea      0.7482 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6678 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.4572 ;
        AntennaPartialMetalArea      0.7115 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5814 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFSHQX4
MACRO DFFSHQX2
    PIN SN
        AntennaGateArea              0.9630 ;
        AntennaPartialMetalArea      4.7713 LAYER met1 ;
        AntennaPartialMetalSideArea  3.7224 LAYER met1 ;
    END SN
    PIN Q
        AntennaPartialMetalArea      1.1814 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7416 LAYER met1 ;
        AntennaDiffArea              1.7967 ;
    END Q
    PIN D
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.7187 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6138 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.6764 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5562 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFSHQX2
MACRO DFFSHQX1
    PIN SN
        AntennaGateArea              0.5688 ;
        AntennaPartialMetalArea      4.3320 LAYER met1 ;
        AntennaPartialMetalSideArea  3.2922 LAYER met1 ;
    END SN
    PIN Q
        AntennaPartialMetalArea      0.8562 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6768 LAYER met1 ;
        AntennaDiffArea              0.9380 ;
    END Q
    PIN D
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.8178 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7650 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2016 ;
        AntennaPartialMetalArea      0.7064 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6174 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFSHQX1
MACRO DFFSXL
    PIN SN
        AntennaGateArea              0.2808 ;
        AntennaPartialMetalArea      2.4847 LAYER met1 ;
        AntennaPartialMetalSideArea  2.3976 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      1.3153 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9666 LAYER met1 ;
        AntennaDiffArea              0.5874 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.7070 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4752 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END Q
    PIN D
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7414 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6750 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7930 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6660 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFSXL
MACRO DFFSX4
    PIN SN
        AntennaGateArea              0.9432 ;
        AntennaPartialMetalArea      3.1977 LAYER met1 ;
        AntennaPartialMetalSideArea  3.1320 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      1.1455 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4590 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8855 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4194 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END Q
    PIN D
        AntennaGateArea              0.1620 ;
        AntennaPartialMetalArea      0.8422 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7092 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7432 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6282 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFSX4
MACRO DFFSX2
    PIN SN
        AntennaGateArea              0.5220 ;
        AntennaPartialMetalArea      2.3342 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2824 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      0.8051 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5904 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.1400 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6624 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Q
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8426 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7722 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.7265 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6012 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFSX2
MACRO DFFSX1
    PIN SN
        AntennaGateArea              0.3348 ;
        AntennaPartialMetalArea      2.3837 LAYER met1 ;
        AntennaPartialMetalSideArea  2.3220 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      1.2994 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9630 LAYER met1 ;
        AntennaDiffArea              0.7732 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6892 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5004 LAYER met1 ;
        AntennaDiffArea              0.8100 ;
    END Q
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7937 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6984 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.7389 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6480 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFSX1
MACRO DFFRHQXL
    PIN RN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9568 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8550 LAYER met1 ;
    END RN
    PIN Q
        AntennaPartialMetalArea      1.0707 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7668 LAYER met1 ;
        AntennaDiffArea              0.9509 ;
    END Q
    PIN D
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.6261 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5598 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6212 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5436 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFRHQXL
MACRO DFFRHQX4
    PIN RN
        AntennaGateArea              0.7380 ;
        AntennaPartialMetalArea      1.0634 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9540 LAYER met1 ;
    END RN
    PIN Q
        AntennaPartialMetalArea      3.0714 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6884 LAYER met1 ;
        AntennaDiffArea              2.8368 ;
    END Q
    PIN D
        AntennaGateArea              0.3348 ;
        AntennaPartialMetalArea      0.8176 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6858 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.4932 ;
        AntennaPartialMetalArea      0.6611 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5544 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFRHQX4
MACRO DFFRHQX2
    PIN RN
        AntennaGateArea              0.4140 ;
        AntennaPartialMetalArea      0.6331 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5490 LAYER met1 ;
    END RN
    PIN Q
        AntennaPartialMetalArea      1.2701 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8730 LAYER met1 ;
        AntennaDiffArea              1.4040 ;
    END Q
    PIN D
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.7906 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7110 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.3060 ;
        AntennaPartialMetalArea      0.6645 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5814 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFRHQX2
MACRO DFFRHQX1
    PIN RN
        AntennaGateArea              0.2628 ;
        AntennaPartialMetalArea      0.8268 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7398 LAYER met1 ;
    END RN
    PIN Q
        AntennaPartialMetalArea      1.0728 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7902 LAYER met1 ;
        AntennaDiffArea              0.9720 ;
    END Q
    PIN D
        AntennaGateArea              0.1332 ;
        AntennaPartialMetalArea      0.6954 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6156 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2160 ;
        AntennaPartialMetalArea      0.7135 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6066 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFRHQX1
MACRO DFFRXL
    PIN RN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6174 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5328 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.2560 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9288 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.5814 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4536 LAYER met1 ;
        AntennaDiffArea              0.6294 ;
    END Q
    PIN D
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.6355 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5922 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7130 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6426 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFRXL
MACRO DFFRX4
    PIN RN
        AntennaGateArea              0.4068 ;
        AntennaPartialMetalArea      1.0354 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9000 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.0640 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5328 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8582 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4410 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END Q
    PIN D
        AntennaGateArea              0.2016 ;
        AntennaPartialMetalArea      0.7845 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7254 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      0.6815 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6030 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFRX4
MACRO DFFRX2
    PIN RN
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      0.7410 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5652 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.9294 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5994 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.1591 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7164 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Q
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6241 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5526 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.7601 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6372 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFRX2
MACRO DFFRX1
    PIN RN
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.6435 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5400 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.3015 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9594 LAYER met1 ;
        AntennaDiffArea              0.7776 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6457 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4716 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7511 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6552 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.6878 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6210 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFRX1
MACRO DFFNSRXL
    PIN SN
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      3.2308 LAYER met1 ;
        AntennaPartialMetalSideArea  2.6496 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.8855 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7506 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.6304 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4680 LAYER met1 ;
        AntennaDiffArea              0.5301 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6060 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4446 LAYER met1 ;
        AntennaDiffArea              0.5674 ;
    END Q
    PIN D
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7259 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6120 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.6470 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5760 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END DFFNSRXL
MACRO DFFNSRX4
    PIN SN
        AntennaGateArea              0.9756 ;
        AntennaPartialMetalArea      4.3592 LAYER met1 ;
        AntennaPartialMetalSideArea  3.5982 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.4428 ;
        AntennaPartialMetalArea      0.7643 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6534 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.9901 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4356 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.0695 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4698 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END Q
    PIN D
        AntennaGateArea              0.2412 ;
        AntennaPartialMetalArea      0.7230 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6462 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.3132 ;
        AntennaPartialMetalArea      0.6451 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5778 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END DFFNSRX4
MACRO DFFNSRX2
    PIN SN
        AntennaGateArea              0.5328 ;
        AntennaPartialMetalArea      3.1839 LAYER met1 ;
        AntennaPartialMetalSideArea  2.6064 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.8444 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7254 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.6796 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5040 LAYER met1 ;
        AntennaDiffArea              1.7040 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.1754 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7776 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Q
    PIN D
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.7086 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6408 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.6726 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6048 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END DFFNSRX2
MACRO DFFNSRX1
    PIN SN
        AntennaGateArea              0.3312 ;
        AntennaPartialMetalArea      3.2276 LAYER met1 ;
        AntennaPartialMetalSideArea  2.6748 LAYER met1 ;
    END SN
    PIN RN
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.8445 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7308 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.9125 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7272 LAYER met1 ;
        AntennaDiffArea              0.7740 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6636 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4734 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN D
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.6944 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6336 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.7118 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6354 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END DFFNSRX1
MACRO DFFNSXL
    PIN SN
        AntennaGateArea              0.2808 ;
        AntennaPartialMetalArea      2.4726 LAYER met1 ;
        AntennaPartialMetalSideArea  2.3886 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      1.2857 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9648 LAYER met1 ;
        AntennaDiffArea              0.5755 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.6870 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4662 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END Q
    PIN D
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.6615 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5796 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6364 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5634 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END DFFNSXL
MACRO DFFNSX4
    PIN SN
        AntennaGateArea              0.9288 ;
        AntennaPartialMetalArea      3.2846 LAYER met1 ;
        AntennaPartialMetalSideArea  3.2202 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      1.4080 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6876 LAYER met1 ;
        AntennaDiffArea              1.5201 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.9924 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5184 LAYER met1 ;
        AntennaDiffArea              1.5201 ;
    END Q
    PIN D
        AntennaGateArea              0.1620 ;
        AntennaPartialMetalArea      0.8116 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6840 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7535 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6426 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END DFFNSX4
MACRO DFFNSX2
    PIN SN
        AntennaGateArea              0.5220 ;
        AntennaPartialMetalArea      2.3718 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2914 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      0.8119 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5652 LAYER met1 ;
        AntennaDiffArea              1.4064 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.2902 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8136 LAYER met1 ;
        AntennaDiffArea              1.5480 ;
    END Q
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9024 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8046 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.8468 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7488 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END DFFNSX2
MACRO DFFNSX1
    PIN SN
        AntennaGateArea              0.3348 ;
        AntennaPartialMetalArea      2.4003 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2734 LAYER met1 ;
    END SN
    PIN QN
        AntennaPartialMetalArea      1.3300 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9972 LAYER met1 ;
        AntennaDiffArea              0.7710 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8116 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4446 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8563 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7596 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.6258 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5580 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END DFFNSX1
MACRO DFFNRXL
    PIN RN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7918 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6894 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.2774 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9630 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.5284 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4338 LAYER met1 ;
        AntennaDiffArea              0.6604 ;
    END Q
    PIN D
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7266 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6192 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7143 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6174 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END DFFNRXL
MACRO DFFNRX4
    PIN RN
        AntennaGateArea              0.3960 ;
        AntennaPartialMetalArea      1.0081 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9270 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.9530 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5310 LAYER met1 ;
        AntennaDiffArea              1.4202 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.8778 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4626 LAYER met1 ;
        AntennaDiffArea              1.4202 ;
    END Q
    PIN D
        AntennaGateArea              0.1980 ;
        AntennaPartialMetalArea      0.6504 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5868 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      0.5945 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5472 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END DFFNRX4
MACRO DFFNRX2
    PIN RN
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      0.7620 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5832 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      0.9294 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5994 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.1770 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7164 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Q
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8339 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7164 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.6798 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6336 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END DFFNRX2
MACRO DFFNRX1
    PIN RN
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.7846 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6822 LAYER met1 ;
    END RN
    PIN QN
        AntennaPartialMetalArea      1.3099 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9828 LAYER met1 ;
        AntennaDiffArea              0.7776 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      0.5708 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4662 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8954 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7614 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1800 ;
        AntennaPartialMetalArea      0.8052 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7092 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END DFFNRX1
MACRO DFFNXL
    PIN QN
        AntennaPartialMetalArea      0.6432 LAYER met1 ;
        AntennaPartialMetalSideArea  0.3978 LAYER met1 ;
        AntennaDiffArea              0.6564 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.1034 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8316 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END Q
    PIN D
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.6710 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6282 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.7294 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6426 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END DFFNXL
MACRO DFFNX4
    PIN QN
        AntennaPartialMetalArea      1.4047 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5166 LAYER met1 ;
        AntennaDiffArea              1.4202 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.0967 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4770 LAYER met1 ;
        AntennaDiffArea              1.4202 ;
    END Q
    PIN D
        AntennaGateArea              0.2988 ;
        AntennaPartialMetalArea      0.7568 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6786 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.4860 ;
        AntennaPartialMetalArea      0.7190 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6480 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END DFFNX4
MACRO DFFNX2
    PIN QN
        AntennaPartialMetalArea      1.0742 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7146 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.1225 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8442 LAYER met1 ;
        AntennaDiffArea              1.0500 ;
    END Q
    PIN D
        AntennaGateArea              0.1620 ;
        AntennaPartialMetalArea      0.7303 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6516 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.6421 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5724 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END DFFNX2
MACRO DFFNX1
    PIN QN
        AntennaPartialMetalArea      0.8220 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4500 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.2313 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9054 LAYER met1 ;
        AntennaDiffArea              0.8040 ;
    END Q
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8833 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7470 LAYER met1 ;
    END D
    PIN CKN
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.8285 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7056 LAYER met1 ;
    END CKN
    PIN GND
    END GND
END DFFNX1
MACRO DFFHQXL
    PIN Q
        AntennaPartialMetalArea      1.0910 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8550 LAYER met1 ;
        AntennaDiffArea              0.6836 ;
    END Q
    PIN D
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.8016 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6822 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.8018 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7470 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFHQXL
MACRO DFFHQX4
    PIN Q
        AntennaPartialMetalArea      1.4154 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7308 LAYER met1 ;
        AntennaDiffArea              1.7640 ;
    END Q
    PIN D
        AntennaGateArea              0.2340 ;
        AntennaPartialMetalArea      0.7814 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7110 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.4140 ;
        AntennaPartialMetalArea      0.6852 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6408 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFHQX4
MACRO DFFHQX2
    PIN Q
        AntennaPartialMetalArea      0.8566 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6354 LAYER met1 ;
        AntennaDiffArea              1.3252 ;
    END Q
    PIN D
        AntennaGateArea              0.1440 ;
        AntennaPartialMetalArea      0.8502 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8064 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2628 ;
        AntennaPartialMetalArea      0.6886 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6210 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFHQX2
MACRO DFFHQX1
    PIN Q
        AntennaPartialMetalArea      1.1132 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8712 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END Q
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8987 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7992 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2016 ;
        AntennaPartialMetalArea      0.7490 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6336 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFHQX1
MACRO DFFXL
    PIN QN
        AntennaPartialMetalArea      0.6432 LAYER met1 ;
        AntennaPartialMetalSideArea  0.3978 LAYER met1 ;
        AntennaDiffArea              0.6564 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.1028 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8280 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END Q
    PIN D
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.8392 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7272 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.8587 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7020 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFXL
MACRO DFFX4
    PIN QN
        AntennaPartialMetalArea      1.4047 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5166 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.0967 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4770 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END Q
    PIN D
        AntennaGateArea              0.2988 ;
        AntennaPartialMetalArea      0.8433 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7236 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.4860 ;
        AntennaPartialMetalArea      0.7333 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6246 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFX4
MACRO DFFX2
    PIN QN
        AntennaPartialMetalArea      1.0742 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7146 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.2297 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8442 LAYER met1 ;
        AntennaDiffArea              1.0500 ;
    END Q
    PIN D
        AntennaGateArea              0.1620 ;
        AntennaPartialMetalArea      0.8137 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7254 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.6672 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5994 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFX2
MACRO DFFX1
    PIN QN
        AntennaPartialMetalArea      0.8153 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5670 LAYER met1 ;
        AntennaDiffArea              0.7860 ;
    END QN
    PIN Q
        AntennaPartialMetalArea      1.4354 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9846 LAYER met1 ;
        AntennaDiffArea              0.8040 ;
    END Q
    PIN D
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.9271 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8208 LAYER met1 ;
    END D
    PIN CK
        AntennaGateArea              0.1908 ;
        AntennaPartialMetalArea      0.7740 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7092 LAYER met1 ;
    END CK
    PIN GND
    END GND
END DFFX1
MACRO CLKINVXL
    PIN Y
        AntennaPartialMetalArea      0.7860 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5868 LAYER met1 ;
        AntennaDiffArea              0.5955 ;
    END Y
    PIN A
        AntennaGateArea              0.1764 ;
        AntennaPartialMetalArea      0.8359 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7326 LAYER met1 ;
    END A
    PIN GND
    END GND
END CLKINVXL
MACRO CLKINVX8
    PIN Y
        AntennaPartialMetalArea      4.3535 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9756 LAYER met1 ;
        AntennaDiffArea              2.4166 ;
    END Y
    PIN A
        AntennaGateArea              1.8572 ;
        AntennaPartialMetalArea      1.4882 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3482 LAYER met1 ;
    END A
    PIN GND
    END GND
END CLKINVX8
MACRO CLKINVX4
    PIN Y
        AntennaPartialMetalArea      1.2316 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6174 LAYER met1 ;
        AntennaDiffArea              1.4273 ;
    END Y
    PIN A
        AntennaGateArea              0.9144 ;
        AntennaPartialMetalArea      0.9943 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8388 LAYER met1 ;
    END A
    PIN GND
    END GND
END CLKINVX4
MACRO CLKINVX3
    PIN Y
        AntennaPartialMetalArea      1.2270 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7218 LAYER met1 ;
        AntennaDiffArea              1.3284 ;
    END Y
    PIN A
        AntennaGateArea              0.6660 ;
        AntennaPartialMetalArea      0.9800 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7758 LAYER met1 ;
    END A
    PIN GND
    END GND
END CLKINVX3
MACRO CLKINVX2
    PIN Y
        AntennaPartialMetalArea      0.9434 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6102 LAYER met1 ;
        AntennaDiffArea              0.8484 ;
    END Y
    PIN A
        AntennaGateArea              0.4392 ;
        AntennaPartialMetalArea      0.8478 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6786 LAYER met1 ;
    END A
    PIN GND
    END GND
END CLKINVX2
MACRO CLKINVX20
    PIN Y
        AntennaPartialMetalArea      16.9800 LAYER met1 ;
        AntennaPartialMetalSideArea  3.3822 LAYER met1 ;
        AntennaDiffArea              12.0277 ;
    END Y
    PIN A
        AntennaGateArea              0.8496 ;
        AntennaPartialMetalArea      1.1308 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8244 LAYER met1 ;
    END A
    PIN GND
    END GND
END CLKINVX20
MACRO CLKINVX1
    PIN Y
        AntennaPartialMetalArea      1.0231 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5454 LAYER met1 ;
        AntennaDiffArea              0.7099 ;
    END Y
    PIN A
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      0.9504 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8064 LAYER met1 ;
    END A
    PIN GND
    END GND
END CLKINVX1
MACRO CLKINVX16
    PIN Y
        AntennaPartialMetalArea      14.5488 LAYER met1 ;
        AntennaPartialMetalSideArea  2.8170 LAYER met1 ;
        AntennaDiffArea              8.5100 ;
    END Y
    PIN A
        AntennaGateArea              0.6732 ;
        AntennaPartialMetalArea      1.0097 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6984 LAYER met1 ;
    END A
    PIN GND
    END GND
END CLKINVX16
MACRO CLKINVX12
    PIN Y
        AntennaPartialMetalArea      12.3230 LAYER met1 ;
        AntennaPartialMetalSideArea  2.5272 LAYER met1 ;
        AntennaDiffArea              6.3946 ;
    END Y
    PIN A
        AntennaGateArea              0.4932 ;
        AntennaPartialMetalArea      0.6809 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6084 LAYER met1 ;
    END A
    PIN GND
    END GND
END CLKINVX12
MACRO CLKBUFXL
    PIN Y
        AntennaPartialMetalArea      0.7954 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5364 LAYER met1 ;
        AntennaDiffArea              0.5940 ;
    END Y
    PIN A
        AntennaGateArea              0.1764 ;
        AntennaPartialMetalArea      0.5776 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5148 LAYER met1 ;
    END A
    PIN GND
    END GND
END CLKBUFXL
MACRO CLKBUFX8
    PIN Y
        AntennaPartialMetalArea      4.4046 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1430 LAYER met1 ;
        AntennaDiffArea              3.1899 ;
    END Y
    PIN A
        AntennaGateArea              0.6192 ;
        AntennaPartialMetalArea      0.9798 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7506 LAYER met1 ;
    END A
    PIN GND
    END GND
END CLKBUFX8
MACRO CLKBUFX4
    PIN Y
        AntennaPartialMetalArea      1.4312 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7020 LAYER met1 ;
        AntennaDiffArea              1.7033 ;
    END Y
    PIN A
        AntennaGateArea              0.2952 ;
        AntennaPartialMetalArea      0.5767 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5166 LAYER met1 ;
    END A
    PIN GND
    END GND
END CLKBUFX4
MACRO CLKBUFX3
    PIN Y
        AntennaPartialMetalArea      1.0428 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6408 LAYER met1 ;
        AntennaDiffArea              1.0734 ;
    END Y
    PIN A
        AntennaGateArea              0.2304 ;
        AntennaPartialMetalArea      0.6022 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5364 LAYER met1 ;
    END A
    PIN GND
    END GND
END CLKBUFX3
MACRO CLKBUFX2
    PIN Y
        AntennaPartialMetalArea      0.7954 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5364 LAYER met1 ;
        AntennaDiffArea              1.3008 ;
    END Y
    PIN A
        AntennaGateArea              0.1944 ;
        AntennaPartialMetalArea      0.5483 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4842 LAYER met1 ;
    END A
    PIN GND
    END GND
END CLKBUFX2
MACRO CLKBUFX20
    PIN Y
        AntennaPartialMetalArea      18.9370 LAYER met1 ;
        AntennaPartialMetalSideArea  3.8052 LAYER met1 ;
        AntennaDiffArea              11.9143 ;
    END Y
    PIN A
        AntennaGateArea              2.4624 ;
        AntennaPartialMetalArea      3.4889 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9638 LAYER met1 ;
    END A
    PIN GND
    END GND
END CLKBUFX20
MACRO CLKBUFX1
    PIN Y
        AntennaPartialMetalArea      0.7984 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5364 LAYER met1 ;
        AntennaDiffArea              0.7084 ;
    END Y
    PIN A
        AntennaGateArea              0.1764 ;
        AntennaPartialMetalArea      0.5483 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4842 LAYER met1 ;
    END A
    PIN GND
    END GND
END CLKBUFX1
MACRO CLKBUFX16
    PIN Y
        AntennaPartialMetalArea      15.6765 LAYER met1 ;
        AntennaPartialMetalSideArea  2.9232 LAYER met1 ;
        AntennaDiffArea              9.6472 ;
    END Y
    PIN A
        AntennaGateArea              2.0124 ;
        AntennaPartialMetalArea      2.9282 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7586 LAYER met1 ;
    END A
    PIN GND
    END GND
END CLKBUFX16
MACRO CLKBUFX12
    PIN Y
        AntennaPartialMetalArea      12.9834 LAYER met1 ;
        AntennaPartialMetalSideArea  2.4714 LAYER met1 ;
        AntennaDiffArea              6.6585 ;
    END Y
    PIN A
        AntennaGateArea              1.5408 ;
        AntennaPartialMetalArea      2.2989 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4454 LAYER met1 ;
    END A
    PIN GND
    END GND
END CLKBUFX12
MACRO BUFXL
    PIN Y
        AntennaPartialMetalArea      0.7878 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5760 LAYER met1 ;
        AntennaDiffArea              0.6172 ;
    END Y
    PIN A
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6586 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5544 LAYER met1 ;
    END A
    PIN GND
    END GND
END BUFXL
MACRO BUFX8
    PIN Y
        AntennaPartialMetalArea      3.2450 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8244 LAYER met1 ;
        AntennaDiffArea              2.8284 ;
    END Y
    PIN A
        AntennaGateArea              0.8820 ;
        AntennaPartialMetalArea      1.0045 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6948 LAYER met1 ;
    END A
    PIN GND
    END GND
END BUFX8
MACRO BUFX4
    PIN Y
        AntennaPartialMetalArea      1.7533 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8154 LAYER met1 ;
        AntennaDiffArea              1.7400 ;
    END Y
    PIN A
        AntennaGateArea              0.4320 ;
        AntennaPartialMetalArea      0.5910 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5148 LAYER met1 ;
    END A
    PIN GND
    END GND
END BUFX4
MACRO BUFX3
    PIN Y
        AntennaPartialMetalArea      1.4976 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7560 LAYER met1 ;
        AntennaDiffArea              1.3108 ;
    END Y
    PIN A
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      0.5707 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5058 LAYER met1 ;
    END A
    PIN GND
    END GND
END BUFX3
MACRO BUFX2
    PIN Y
        AntennaPartialMetalArea      0.8646 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6084 LAYER met1 ;
        AntennaDiffArea              1.6020 ;
    END Y
    PIN A
        AntennaGateArea              0.2160 ;
        AntennaPartialMetalArea      0.5898 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5220 LAYER met1 ;
    END A
    PIN GND
    END GND
END BUFX2
MACRO BUFX20
    PIN Y
        AntennaPartialMetalArea      11.3606 LAYER met1 ;
        AntennaPartialMetalSideArea  2.6118 LAYER met1 ;
        AntennaDiffArea              7.8122 ;
    END Y
    PIN A
        AntennaGateArea              2.2032 ;
        AntennaPartialMetalArea      2.6218 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6650 LAYER met1 ;
    END A
    PIN GND
    END GND
END BUFX20
MACRO BUFX1
    PIN Y
        AntennaPartialMetalArea      0.6815 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5004 LAYER met1 ;
        AntennaDiffArea              0.8250 ;
    END Y
    PIN A
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6374 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5634 LAYER met1 ;
    END A
    PIN GND
    END GND
END BUFX1
MACRO BUFX16
    PIN Y
        AntennaPartialMetalArea      9.3900 LAYER met1 ;
        AntennaPartialMetalSideArea  2.1420 LAYER met1 ;
        AntennaDiffArea              6.3596 ;
    END Y
    PIN A
        AntennaGateArea              1.7496 ;
        AntennaPartialMetalArea      2.0904 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2744 LAYER met1 ;
    END A
    PIN GND
    END GND
END BUFX16
MACRO BUFX12
    PIN Y
        AntennaPartialMetalArea      6.5537 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4562 LAYER met1 ;
        AntennaDiffArea              4.2426 ;
    END Y
    PIN A
        AntennaGateArea              1.3032 ;
        AntennaPartialMetalArea      1.3807 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9684 LAYER met1 ;
    END A
    PIN GND
    END GND
END BUFX12
MACRO AOI33XL
    PIN Y
        AntennaPartialMetalArea      1.8860 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3878 LAYER met1 ;
        AntennaDiffArea              1.3398 ;
    END Y
    PIN B2
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.8727 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6804 LAYER met1 ;
    END B2
    PIN B1
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.7602 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6732 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.6884 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6156 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.7252 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6534 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.7065 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6282 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.8274 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7236 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI33XL
MACRO AOI33X4
    PIN Y
        AntennaPartialMetalArea      0.8955 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4482 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END Y
    PIN B2
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.9007 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7596 LAYER met1 ;
    END B2
    PIN B1
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.8146 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7362 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.8282 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7560 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.8732 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8028 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.8803 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8226 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.8212 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7686 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI33X4
MACRO AOI33X2
    PIN Y
        AntennaPartialMetalArea      3.8468 LAYER met1 ;
        AntennaPartialMetalSideArea  2.5344 LAYER met1 ;
        AntennaDiffArea              2.7495 ;
    END Y
    PIN B2
        AntennaGateArea              0.7920 ;
        AntennaPartialMetalArea      2.2536 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8684 LAYER met1 ;
    END B2
    PIN B1
        AntennaGateArea              0.7920 ;
        AntennaPartialMetalArea      1.8339 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5804 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.7920 ;
        AntennaPartialMetalArea      1.0959 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9954 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.7920 ;
        AntennaPartialMetalArea      2.2638 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8792 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.7920 ;
        AntennaPartialMetalArea      1.7991 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6740 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.7920 ;
        AntennaPartialMetalArea      1.2816 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0188 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI33X2
MACRO AOI33X1
    PIN Y
        AntennaPartialMetalArea      1.8981 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3824 LAYER met1 ;
        AntennaDiffArea              1.9248 ;
    END Y
    PIN B2
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.9541 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7704 LAYER met1 ;
    END B2
    PIN B1
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.7976 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7200 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.6774 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6030 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.6948 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6372 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.6939 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6156 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.8220 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7164 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI33X1
MACRO AOI32XL
    PIN Y
        AntennaPartialMetalArea      1.5901 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1268 LAYER met1 ;
        AntennaDiffArea              0.8900 ;
    END Y
    PIN B1
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.8397 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7848 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7871 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7272 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.9151 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7740 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.9114 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7992 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.8399 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7722 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI32XL
MACRO AOI32X4
    PIN Y
        AntennaPartialMetalArea      0.8485 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4680 LAYER met1 ;
        AntennaDiffArea              1.4142 ;
    END Y
    PIN B1
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      0.8609 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8118 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      0.8208 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7254 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.9007 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7596 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.8146 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7362 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.8249 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7578 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI32X4
MACRO AOI32X2
    PIN Y
        AntennaPartialMetalArea      2.8352 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8900 LAYER met1 ;
        AntennaDiffArea              2.1556 ;
    END Y
    PIN B1
        AntennaGateArea              0.7344 ;
        AntennaPartialMetalArea      1.7184 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4436 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.7344 ;
        AntennaPartialMetalArea      1.1022 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9936 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.7920 ;
        AntennaPartialMetalArea      2.1340 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8306 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.7920 ;
        AntennaPartialMetalArea      1.7713 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5282 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.7920 ;
        AntennaPartialMetalArea      1.0980 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0332 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI32X2
MACRO AOI32X1
    PIN Y
        AntennaPartialMetalArea      1.4284 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0638 LAYER met1 ;
        AntennaDiffArea              1.2272 ;
    END Y
    PIN B1
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7551 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7002 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7025 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6426 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.8206 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6750 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.8510 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7128 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.7448 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6714 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI32X1
MACRO AOI31XL
    PIN Y
        AntennaPartialMetalArea      1.0340 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7776 LAYER met1 ;
        AntennaDiffArea              0.8166 ;
    END Y
    PIN B0
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      0.7484 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7074 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.7976 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7002 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.7733 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6894 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2700 ;
        AntennaPartialMetalArea      0.8088 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7254 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI31XL
MACRO AOI31X4
    PIN Y
        AntennaPartialMetalArea      1.5166 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7668 LAYER met1 ;
        AntennaDiffArea              1.4526 ;
    END Y
    PIN B0
        AntennaGateArea              0.2052 ;
        AntennaPartialMetalArea      0.7088 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6048 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.8343 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7272 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.8674 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7002 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2448 ;
        AntennaPartialMetalArea      0.6312 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5814 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI31X4
MACRO AOI31X2
    PIN Y
        AntennaPartialMetalArea      2.0970 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4706 LAYER met1 ;
        AntennaDiffArea              1.7541 ;
    END Y
    PIN B0
        AntennaGateArea              0.6624 ;
        AntennaPartialMetalArea      1.0388 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8874 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.7920 ;
        AntennaPartialMetalArea      1.3909 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1790 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.7920 ;
        AntennaPartialMetalArea      1.6587 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4400 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.7920 ;
        AntennaPartialMetalArea      2.1260 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8180 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI31X2
MACRO AOI31X1
    PIN Y
        AntennaPartialMetalArea      1.2328 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8982 LAYER met1 ;
        AntennaDiffArea              1.0909 ;
    END Y
    PIN B0
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      0.8222 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7776 LAYER met1 ;
    END B0
    PIN A2
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.8732 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7038 LAYER met1 ;
    END A2
    PIN A1
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.8734 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6786 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.3888 ;
        AntennaPartialMetalArea      0.8317 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7038 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI31X1
MACRO AOI2BB2XL
    PIN Y
        AntennaPartialMetalArea      0.9165 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7092 LAYER met1 ;
        AntennaDiffArea              0.7677 ;
    END Y
    PIN B1
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7963 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7092 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.8608 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7290 LAYER met1 ;
    END B0
    PIN A1N
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.8854 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7776 LAYER met1 ;
    END A1N
    PIN A0N
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.8551 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7722 LAYER met1 ;
    END A0N
    PIN GND
    END GND
END AOI2BB2XL
MACRO AOI2BB2X4
    PIN Y
        AntennaPartialMetalArea      4.2856 LAYER met1 ;
        AntennaPartialMetalSideArea  2.4840 LAYER met1 ;
        AntennaDiffArea              3.4904 ;
    END Y
    PIN B1
        AntennaGateArea              1.4562 ;
        AntennaPartialMetalArea      3.1265 LAYER met1 ;
        AntennaPartialMetalSideArea  2.4678 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              1.4562 ;
        AntennaPartialMetalArea      2.2232 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6848 LAYER met1 ;
    END B0
    PIN A1N
        AntennaGateArea              0.6048 ;
        AntennaPartialMetalArea      1.9094 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5732 LAYER met1 ;
    END A1N
    PIN A0N
        AntennaGateArea              0.6048 ;
        AntennaPartialMetalArea      0.9966 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8208 LAYER met1 ;
    END A0N
    PIN GND
    END GND
END AOI2BB2X4
MACRO AOI2BB2X2
    PIN Y
        AntennaPartialMetalArea      1.9776 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4382 LAYER met1 ;
        AntennaDiffArea              1.6860 ;
    END Y
    PIN B1
        AntennaGateArea              0.7344 ;
        AntennaPartialMetalArea      1.9295 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6506 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.7344 ;
        AntennaPartialMetalArea      2.1753 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7964 LAYER met1 ;
    END B0
    PIN A1N
        AntennaGateArea              0.3132 ;
        AntennaPartialMetalArea      0.6575 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5958 LAYER met1 ;
    END A1N
    PIN A0N
        AntennaGateArea              0.3132 ;
        AntennaPartialMetalArea      0.7930 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6570 LAYER met1 ;
    END A0N
    PIN GND
    END GND
END AOI2BB2X2
MACRO AOI2BB2X1
    PIN Y
        AntennaPartialMetalArea      1.2848 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9702 LAYER met1 ;
        AntennaDiffArea              0.9195 ;
    END Y
    PIN B1
        AntennaGateArea              0.3672 ;
        AntennaPartialMetalArea      0.7760 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7092 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.3672 ;
        AntennaPartialMetalArea      0.7230 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6750 LAYER met1 ;
    END B0
    PIN A1N
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.7742 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6966 LAYER met1 ;
    END A1N
    PIN A0N
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.7739 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7074 LAYER met1 ;
    END A0N
    PIN GND
    END GND
END AOI2BB2X1
MACRO AOI2BB1XL
    PIN Y
        AntennaPartialMetalArea      0.8794 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6876 LAYER met1 ;
        AntennaDiffArea              0.7036 ;
    END Y
    PIN B0
        AntennaGateArea              0.2340 ;
        AntennaPartialMetalArea      0.8462 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7200 LAYER met1 ;
    END B0
    PIN A1N
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.7489 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6642 LAYER met1 ;
    END A1N
    PIN A0N
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.9634 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8550 LAYER met1 ;
    END A0N
    PIN GND
    END GND
END AOI2BB1XL
MACRO AOI2BB1X4
    PIN Y
        AntennaPartialMetalArea      3.4080 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7424 LAYER met1 ;
        AntennaDiffArea              2.7358 ;
    END Y
    PIN B0
        AntennaGateArea              1.3290 ;
        AntennaPartialMetalArea      1.4645 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3968 LAYER met1 ;
    END B0
    PIN A1N
        AntennaGateArea              0.6156 ;
        AntennaPartialMetalArea      2.0774 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6884 LAYER met1 ;
    END A1N
    PIN A0N
        AntennaGateArea              0.6156 ;
        AntennaPartialMetalArea      0.9253 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7758 LAYER met1 ;
    END A0N
    PIN GND
    END GND
END AOI2BB1X4
MACRO AOI2BB1X2
    PIN Y
        AntennaPartialMetalArea      1.6084 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1538 LAYER met1 ;
        AntennaDiffArea              1.3920 ;
    END Y
    PIN B0
        AntennaGateArea              0.6480 ;
        AntennaPartialMetalArea      1.3596 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1232 LAYER met1 ;
    END B0
    PIN A1N
        AntennaGateArea              0.3132 ;
        AntennaPartialMetalArea      0.7368 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6534 LAYER met1 ;
    END A1N
    PIN A0N
        AntennaGateArea              0.3132 ;
        AntennaPartialMetalArea      0.7603 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6156 LAYER met1 ;
    END A0N
    PIN GND
    END GND
END AOI2BB1X2
MACRO AOI2BB1X1
    PIN Y
        AntennaPartialMetalArea      0.9809 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7758 LAYER met1 ;
        AntennaDiffArea              0.9527 ;
    END Y
    PIN B0
        AntennaGateArea              0.3168 ;
        AntennaPartialMetalArea      0.8038 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7074 LAYER met1 ;
    END B0
    PIN A1N
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      0.7331 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6552 LAYER met1 ;
    END A1N
    PIN A0N
        AntennaGateArea              0.1548 ;
        AntennaPartialMetalArea      1.0105 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8946 LAYER met1 ;
    END A0N
    PIN GND
    END GND
END AOI2BB1X1
MACRO AOI22XL
    PIN Y
        AntennaPartialMetalArea      1.3946 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0476 LAYER met1 ;
        AntennaDiffArea              0.8120 ;
    END Y
    PIN B1
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7920 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6696 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7654 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6390 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7560 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6822 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7897 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6606 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI22XL
MACRO AOI22X4
    PIN Y
        AntennaPartialMetalArea      7.4932 LAYER met1 ;
        AntennaPartialMetalSideArea  3.1842 LAYER met1 ;
        AntennaDiffArea              5.4740 ;
    END Y
    PIN B1
        AntennaGateArea              1.4610 ;
        AntennaPartialMetalArea      2.4619 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8540 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              1.4610 ;
        AntennaPartialMetalArea      2.4601 LAYER met1 ;
        AntennaPartialMetalSideArea  2.0700 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              1.4610 ;
        AntennaPartialMetalArea      2.2425 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8972 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              1.4610 ;
        AntennaPartialMetalArea      2.5022 LAYER met1 ;
        AntennaPartialMetalSideArea  1.9872 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI22X4
MACRO AOI22X2
    PIN Y
        AntennaPartialMetalArea      2.2188 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6614 LAYER met1 ;
        AntennaDiffArea              2.1079 ;
    END Y
    PIN B1
        AntennaGateArea              0.7344 ;
        AntennaPartialMetalArea      2.0914 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4760 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.7344 ;
        AntennaPartialMetalArea      1.4672 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1304 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.7344 ;
        AntennaPartialMetalArea      1.7131 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4418 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.7344 ;
        AntennaPartialMetalArea      1.2163 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0098 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI22X2
MACRO AOI22X1
    PIN Y
        AntennaPartialMetalArea      1.4022 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0584 LAYER met1 ;
        AntennaDiffArea              1.1600 ;
    END Y
    PIN B1
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7278 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6282 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7991 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6444 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7788 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6840 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7388 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6930 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI22X1
MACRO AOI222XL
    PIN Y
        AntennaPartialMetalArea      2.0696 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5930 LAYER met1 ;
        AntennaDiffArea              1.1689 ;
    END Y
    PIN C1
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      0.7480 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6678 LAYER met1 ;
    END C1
    PIN C0
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      0.7786 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6966 LAYER met1 ;
    END C0
    PIN B1
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      0.9224 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7434 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      0.7668 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6948 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      0.6770 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6336 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      0.6899 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6138 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI222XL
MACRO AOI222X4
    PIN Y
        AntennaPartialMetalArea      1.0456 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6282 LAYER met1 ;
        AntennaDiffArea              1.6872 ;
    END Y
    PIN C1
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.7238 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6318 LAYER met1 ;
    END C1
    PIN C0
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.7477 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6246 LAYER met1 ;
    END C0
    PIN B1
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.8069 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6588 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.6154 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5454 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.8045 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6840 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.7274 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6714 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI222X4
MACRO AOI222X2
    PIN Y
        AntennaPartialMetalArea      3.3502 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2698 LAYER met1 ;
        AntennaDiffArea              2.6242 ;
    END Y
    PIN C1
        AntennaGateArea              0.8064 ;
        AntennaPartialMetalArea      1.4882 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2672 LAYER met1 ;
    END C1
    PIN C0
        AntennaGateArea              0.8064 ;
        AntennaPartialMetalArea      1.0088 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8640 LAYER met1 ;
    END C0
    PIN B1
        AntennaGateArea              0.8064 ;
        AntennaPartialMetalArea      1.7926 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4976 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.8064 ;
        AntennaPartialMetalArea      1.0452 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9828 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.8064 ;
        AntennaPartialMetalArea      1.6990 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4994 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.8064 ;
        AntennaPartialMetalArea      1.0880 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9954 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI222X2
MACRO AOI222X1
    PIN Y
        AntennaPartialMetalArea      2.4217 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7964 LAYER met1 ;
        AntennaDiffArea              1.6481 ;
    END Y
    PIN C1
        AntennaGateArea              0.4032 ;
        AntennaPartialMetalArea      0.6562 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5796 LAYER met1 ;
    END C1
    PIN C0
        AntennaGateArea              0.4032 ;
        AntennaPartialMetalArea      0.6688 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6156 LAYER met1 ;
    END C0
    PIN B1
        AntennaGateArea              0.4032 ;
        AntennaPartialMetalArea      0.7214 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6804 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.4032 ;
        AntennaPartialMetalArea      0.7875 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7182 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.4032 ;
        AntennaPartialMetalArea      1.0396 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7884 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.4032 ;
        AntennaPartialMetalArea      0.8553 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7776 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI222X1
MACRO AOI221XL
    PIN Y
        AntennaPartialMetalArea      1.3598 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0080 LAYER met1 ;
        AntennaDiffArea              1.1295 ;
    END Y
    PIN C0
        AntennaGateArea              0.2628 ;
        AntennaPartialMetalArea      0.7389 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6786 LAYER met1 ;
    END C0
    PIN B1
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      0.7902 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7344 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      0.8237 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7236 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      0.8135 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7650 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2880 ;
        AntennaPartialMetalArea      0.7657 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7218 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI221XL
MACRO AOI221X4
    PIN Y
        AntennaPartialMetalArea      1.2987 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6984 LAYER met1 ;
        AntennaDiffArea              1.7400 ;
    END Y
    PIN C0
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      0.8322 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7596 LAYER met1 ;
    END C0
    PIN B1
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.7442 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6912 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.7467 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6840 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.8002 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7236 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.8276 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7506 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI221X4
MACRO AOI221X2
    PIN Y
        AntennaPartialMetalArea      2.4605 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8108 LAYER met1 ;
        AntennaDiffArea              2.1036 ;
    END Y
    PIN C0
        AntennaGateArea              0.7332 ;
        AntennaPartialMetalArea      1.3060 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0170 LAYER met1 ;
    END C0
    PIN B1
        AntennaGateArea              0.8052 ;
        AntennaPartialMetalArea      1.5996 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3968 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.8052 ;
        AntennaPartialMetalArea      1.3688 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1070 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.8052 ;
        AntennaPartialMetalArea      1.8117 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5570 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.8052 ;
        AntennaPartialMetalArea      1.2361 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0116 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI221X2
MACRO AOI221X1
    PIN Y
        AntennaPartialMetalArea      1.4125 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0314 LAYER met1 ;
        AntennaDiffArea              1.3242 ;
    END Y
    PIN C0
        AntennaGateArea              0.3666 ;
        AntennaPartialMetalArea      0.7616 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6966 LAYER met1 ;
    END C0
    PIN B1
        AntennaGateArea              0.4026 ;
        AntennaPartialMetalArea      0.7280 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6462 LAYER met1 ;
    END B1
    PIN B0
        AntennaGateArea              0.4026 ;
        AntennaPartialMetalArea      0.7178 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6552 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.4026 ;
        AntennaPartialMetalArea      0.8291 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7758 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.4026 ;
        AntennaPartialMetalArea      0.8136 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7182 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI221X1
MACRO AOI21XL
    PIN Y
        AntennaPartialMetalArea      1.1636 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8388 LAYER met1 ;
        AntennaDiffArea              0.8083 ;
    END Y
    PIN B0
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      0.8260 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7020 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.9324 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7848 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7518 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6786 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI21XL
MACRO AOI21X4
    PIN Y
        AntennaPartialMetalArea      4.7226 LAYER met1 ;
        AntennaPartialMetalSideArea  2.2482 LAYER met1 ;
        AntennaDiffArea              3.3352 ;
    END Y
    PIN B0
        AntennaGateArea              1.3250 ;
        AntennaPartialMetalArea      1.9480 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3482 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              1.4610 ;
        AntennaPartialMetalArea      2.0769 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6992 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              1.4610 ;
        AntennaPartialMetalArea      2.3703 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8432 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI21X4
MACRO AOI21X2
    PIN Y
        AntennaPartialMetalArea      1.6955 LAYER met1 ;
        AntennaPartialMetalSideArea  1.2618 LAYER met1 ;
        AntennaDiffArea              1.6348 ;
    END Y
    PIN B0
        AntennaGateArea              0.6696 ;
        AntennaPartialMetalArea      0.8744 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7686 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.7344 ;
        AntennaPartialMetalArea      1.0483 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9738 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.7344 ;
        AntennaPartialMetalArea      1.7637 LAYER met1 ;
        AntennaPartialMetalSideArea  1.4904 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI21X2
MACRO AOI21X1
    PIN Y
        AntennaPartialMetalArea      1.1662 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8244 LAYER met1 ;
        AntennaDiffArea              1.1160 ;
    END Y
    PIN B0
        AntennaGateArea              0.3240 ;
        AntennaPartialMetalArea      0.6292 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5364 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7233 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5760 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7620 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6480 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI21X1
MACRO AOI211XL
    PIN Y
        AntennaPartialMetalArea      1.2321 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9666 LAYER met1 ;
        AntennaDiffArea              1.2157 ;
    END Y
    PIN C0
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.7226 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6372 LAYER met1 ;
    END C0
    PIN B0
        AntennaGateArea              0.2520 ;
        AntennaPartialMetalArea      0.6374 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5706 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.7276 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6606 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.9000 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7902 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI211XL
MACRO AOI211X4
    PIN Y
        AntennaPartialMetalArea      1.3057 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6480 LAYER met1 ;
        AntennaDiffArea              1.5922 ;
    END Y
    PIN C0
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      0.7058 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6282 LAYER met1 ;
    END C0
    PIN B0
        AntennaGateArea              0.2268 ;
        AntennaPartialMetalArea      0.9828 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8406 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.6958 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6192 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.2484 ;
        AntennaPartialMetalArea      0.7901 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6804 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI211X4
MACRO AOI211X2
    PIN Y
        AntennaPartialMetalArea      2.4872 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7172 LAYER met1 ;
        AntennaDiffArea              2.8152 ;
    END Y
    PIN C0
        AntennaGateArea              0.7200 ;
        AntennaPartialMetalArea      1.4078 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1646 LAYER met1 ;
    END C0
    PIN B0
        AntennaGateArea              0.7200 ;
        AntennaPartialMetalArea      0.7914 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6894 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.8084 ;
        AntennaPartialMetalArea      1.1167 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0368 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.8068 ;
        AntennaPartialMetalArea      1.6150 LAYER met1 ;
        AntennaPartialMetalSideArea  1.3320 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI211X2
MACRO AOI211X1
    PIN Y
        AntennaPartialMetalArea      1.8742 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1016 LAYER met1 ;
        AntennaDiffArea              1.4240 ;
    END Y
    PIN C0
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7885 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6822 LAYER met1 ;
    END C0
    PIN B0
        AntennaGateArea              0.3600 ;
        AntennaPartialMetalArea      0.7628 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6156 LAYER met1 ;
    END B0
    PIN A1
        AntennaGateArea              0.3960 ;
        AntennaPartialMetalArea      0.7817 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6426 LAYER met1 ;
    END A1
    PIN A0
        AntennaGateArea              0.3960 ;
        AntennaPartialMetalArea      0.7644 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6660 LAYER met1 ;
    END A0
    PIN GND
    END GND
END AOI211X1
MACRO ANTENNA
    CLASS CORE ANTENNACELL ;
    PIN A
        AntennaPartialMetalArea      0.4154 LAYER met1 ;
        AntennaPartialMetalSideArea  0.2322 LAYER met1 ;
        AntennaDiffArea              1.1128 ;
    END A
    PIN GND
    END GND
END ANTENNA
MACRO AND4XL
    PIN Y
        AntennaPartialMetalArea      0.6804 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5508 LAYER met1 ;
        AntennaDiffArea              0.5899 ;
    END Y
    PIN D
        AntennaGateArea              0.1584 ;
        AntennaPartialMetalArea      0.9226 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7704 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.1584 ;
        AntennaPartialMetalArea      0.8220 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7092 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.1584 ;
        AntennaPartialMetalArea      0.8166 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7002 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.1584 ;
        AntennaPartialMetalArea      1.0458 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9774 LAYER met1 ;
    END A
    PIN GND
    END GND
END AND4XL
MACRO AND4X4
    PIN Y
        AntennaPartialMetalArea      1.1936 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7452 LAYER met1 ;
        AntennaDiffArea              1.6072 ;
    END Y
    PIN D
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.8626 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6750 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.7626 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6714 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.7302 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6552 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.7972 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6984 LAYER met1 ;
    END A
    PIN GND
    END GND
END AND4X4
MACRO AND4X2
    PIN Y
        AntennaPartialMetalArea      1.0712 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7110 LAYER met1 ;
        AntennaDiffArea              1.3980 ;
    END Y
    PIN D
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.9229 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8010 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.8319 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7200 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.8426 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7704 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.2772 ;
        AntennaPartialMetalArea      0.9261 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7866 LAYER met1 ;
    END A
    PIN GND
    END GND
END AND4X2
MACRO AND4X1
    PIN Y
        AntennaPartialMetalArea      0.7548 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5886 LAYER met1 ;
        AntennaDiffArea              0.7687 ;
    END Y
    PIN D
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.9191 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7704 LAYER met1 ;
    END D
    PIN C
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.8290 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6984 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.7788 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6822 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.1368 ;
        AntennaPartialMetalArea      0.9918 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9234 LAYER met1 ;
    END A
    PIN GND
    END GND
END AND4X1
MACRO AND3XL
    PIN Y
        AntennaPartialMetalArea      0.8567 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6228 LAYER met1 ;
        AntennaDiffArea              0.5913 ;
    END Y
    PIN C
        AntennaGateArea              0.1512 ;
        AntennaPartialMetalArea      0.8196 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7524 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.1512 ;
        AntennaPartialMetalArea      1.0524 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9810 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.1512 ;
        AntennaPartialMetalArea      1.1153 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0512 LAYER met1 ;
    END A
    PIN GND
    END GND
END AND3XL
MACRO AND3X4
    PIN Y
        AntennaPartialMetalArea      1.4802 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7164 LAYER met1 ;
        AntennaDiffArea              1.7400 ;
    END Y
    PIN C
        AntennaGateArea              0.5220 ;
        AntennaPartialMetalArea      0.6008 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5382 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.5220 ;
        AntennaPartialMetalArea      0.6437 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5652 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5220 ;
        AntennaPartialMetalArea      0.8511 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7020 LAYER met1 ;
    END A
    PIN GND
    END GND
END AND3X4
MACRO AND3X2
    PIN Y
        AntennaPartialMetalArea      0.9600 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6516 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Y
    PIN C
        AntennaGateArea              0.2664 ;
        AntennaPartialMetalArea      0.7882 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6858 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.2664 ;
        AntennaPartialMetalArea      0.7550 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6228 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.2664 ;
        AntennaPartialMetalArea      0.7454 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6570 LAYER met1 ;
    END A
    PIN GND
    END GND
END AND3X2
MACRO AND3X1
    PIN Y
        AntennaPartialMetalArea      0.9523 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7362 LAYER met1 ;
        AntennaDiffArea              0.7764 ;
    END Y
    PIN C
        AntennaGateArea              0.1332 ;
        AntennaPartialMetalArea      0.9066 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8208 LAYER met1 ;
    END C
    PIN B
        AntennaGateArea              0.1332 ;
        AntennaPartialMetalArea      1.1094 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0314 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.1332 ;
        AntennaPartialMetalArea      1.1336 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0620 LAYER met1 ;
    END A
    PIN GND
    END GND
END AND3X1
MACRO AND2XL
    PIN Y
        AntennaPartialMetalArea      0.5578 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4608 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END Y
    PIN B
        AntennaGateArea              0.1332 ;
        AntennaPartialMetalArea      0.6689 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5832 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.1332 ;
        AntennaPartialMetalArea      0.8914 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8262 LAYER met1 ;
    END A
    PIN GND
    END GND
END AND2XL
MACRO AND2X4
    PIN Y
        AntennaPartialMetalArea      1.2627 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6534 LAYER met1 ;
        AntennaDiffArea              1.4481 ;
    END Y
    PIN B
        AntennaGateArea              0.4392 ;
        AntennaPartialMetalArea      0.7820 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6840 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.4392 ;
        AntennaPartialMetalArea      0.6776 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6084 LAYER met1 ;
    END A
    PIN GND
    END GND
END AND2X4
MACRO AND2X2
    PIN Y
        AntennaPartialMetalArea      1.3662 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6660 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END Y
    PIN B
        AntennaGateArea              0.2376 ;
        AntennaPartialMetalArea      0.7566 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6552 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.2376 ;
        AntennaPartialMetalArea      0.8369 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6822 LAYER met1 ;
    END A
    PIN GND
    END GND
END AND2X2
MACRO AND2X1
    PIN Y
        AntennaPartialMetalArea      0.5724 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4716 LAYER met1 ;
        AntennaDiffArea              0.7477 ;
    END Y
    PIN B
        AntennaGateArea              0.1224 ;
        AntennaPartialMetalArea      0.6728 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5868 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.1224 ;
        AntennaPartialMetalArea      0.9180 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8280 LAYER met1 ;
    END A
    PIN GND
    END GND
END AND2X1
MACRO ADDHXL
    PIN S
        AntennaPartialMetalArea      1.0398 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8010 LAYER met1 ;
        AntennaDiffArea              1.2260 ;
    END S
    PIN CO
        AntennaPartialMetalArea      0.6316 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4734 LAYER met1 ;
        AntennaDiffArea              0.6214 ;
    END CO
    PIN B
        AntennaGateArea              0.5220 ;
        AntennaPartialMetalArea      3.9728 LAYER met1 ;
        AntennaPartialMetalSideArea  3.1266 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.3312 ;
        AntennaPartialMetalArea      1.4028 LAYER met1 ;
        AntennaPartialMetalSideArea  1.1070 LAYER met1 ;
    END A
    PIN GND
    END GND
END ADDHXL
MACRO ADDHX4
    PIN S
        AntennaPartialMetalArea      5.4490 LAYER met1 ;
        AntennaPartialMetalSideArea  2.5920 LAYER met1 ;
        AntennaDiffArea              7.3085 ;
    END S
    PIN CO
        AntennaPartialMetalArea      1.8814 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8874 LAYER met1 ;
        AntennaDiffArea              1.4652 ;
    END CO
    PIN B
        AntennaGateArea              3.5640 ;
        AntennaPartialMetalArea      4.9107 LAYER met1 ;
        AntennaPartialMetalSideArea  3.8394 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              3.5604 ;
        AntennaPartialMetalArea      4.1802 LAYER met1 ;
        AntennaPartialMetalSideArea  2.9610 LAYER met1 ;
    END A
    PIN GND
    END GND
END ADDHX4
MACRO ADDHX2
    PIN S
        AntennaPartialMetalArea      2.1083 LAYER met1 ;
        AntennaPartialMetalSideArea  1.5948 LAYER met1 ;
        AntennaDiffArea              3.9951 ;
    END S
    PIN CO
        AntennaPartialMetalArea      0.7948 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4950 LAYER met1 ;
        AntennaDiffArea              1.2455 ;
    END CO
    PIN B
        AntennaGateArea              1.7748 ;
        AntennaPartialMetalArea      2.8080 LAYER met1 ;
        AntennaPartialMetalSideArea  2.3562 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              1.8000 ;
        AntennaPartialMetalArea      2.3276 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7046 LAYER met1 ;
    END A
    PIN GND
    END GND
END ADDHX2
MACRO ADDHX1
    PIN S
        AntennaPartialMetalArea      1.0398 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8010 LAYER met1 ;
        AntennaDiffArea              2.3880 ;
    END S
    PIN CO
        AntennaPartialMetalArea      0.7970 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5850 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END CO
    PIN B
        AntennaGateArea              0.8784 ;
        AntennaPartialMetalArea      4.3095 LAYER met1 ;
        AntennaPartialMetalSideArea  3.4434 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.8784 ;
        AntennaPartialMetalArea      1.4427 LAYER met1 ;
        AntennaPartialMetalSideArea  1.0926 LAYER met1 ;
    END A
    PIN GND
    END GND
END ADDHX1
MACRO ADDFHXL
    PIN S
        AntennaPartialMetalArea      0.8178 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5706 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END S
    PIN CO
        AntennaPartialMetalArea      0.6817 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5112 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END CO
    PIN CI
        AntennaGateArea              0.1296 ;
        AntennaPartialMetalArea      0.6980 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5886 LAYER met1 ;
    END CI
    PIN B
        AntennaGateArea              0.6336 ;
        AntennaPartialMetalArea      2.9788 LAYER met1 ;
        AntennaPartialMetalSideArea  2.8188 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.2592 ;
        AntennaPartialMetalArea      0.8768 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7974 LAYER met1 ;
    END A
    PIN GND
    END GND
END ADDFHXL
MACRO ADDFHX4
    PIN S
        AntennaPartialMetalArea      0.8440 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4338 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END S
    PIN CO
        AntennaPartialMetalArea      0.9410 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4734 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END CO
    PIN CI
        AntennaGateArea              0.6048 ;
        AntennaPartialMetalArea      1.2508 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9540 LAYER met1 ;
    END CI
    PIN B
        AntennaGateArea              2.3256 ;
        AntennaPartialMetalArea      4.7575 LAYER met1 ;
        AntennaPartialMetalSideArea  4.0788 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.9684 ;
        AntennaPartialMetalArea      1.1936 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9306 LAYER met1 ;
    END A
    PIN GND
    END GND
END ADDFHX4
MACRO ADDFHX2
    PIN S
        AntennaPartialMetalArea      1.1412 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6966 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END S
    PIN CO
        AntennaPartialMetalArea      0.6614 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4932 LAYER met1 ;
        AntennaDiffArea              1.5030 ;
    END CO
    PIN CI
        AntennaGateArea              0.6048 ;
        AntennaPartialMetalArea      1.2851 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9378 LAYER met1 ;
    END CI
    PIN B
        AntennaGateArea              2.3112 ;
        AntennaPartialMetalArea      4.8273 LAYER met1 ;
        AntennaPartialMetalSideArea  4.0986 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.9684 ;
        AntennaPartialMetalArea      1.1696 LAYER met1 ;
        AntennaPartialMetalSideArea  0.9216 LAYER met1 ;
    END A
    PIN GND
    END GND
END ADDFHX2
MACRO ADDFHX1
    PIN S
        AntennaPartialMetalArea      0.8202 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6066 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END S
    PIN CO
        AntennaPartialMetalArea      0.7388 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5130 LAYER met1 ;
        AntennaDiffArea              0.7860 ;
    END CO
    PIN CI
        AntennaGateArea              0.2988 ;
        AntennaPartialMetalArea      0.7207 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5958 LAYER met1 ;
    END CI
    PIN B
        AntennaGateArea              1.1700 ;
        AntennaPartialMetalArea      3.6177 LAYER met1 ;
        AntennaPartialMetalSideArea  3.1284 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.4788 ;
        AntennaPartialMetalArea      0.9360 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7524 LAYER met1 ;
    END A
    PIN GND
    END GND
END ADDFHX1
MACRO ADDFXL
    PIN S
        AntennaPartialMetalArea      0.6570 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4770 LAYER met1 ;
        AntennaDiffArea              0.5825 ;
    END S
    PIN CO
        AntennaPartialMetalArea      0.6478 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4338 LAYER met1 ;
        AntennaDiffArea              0.5810 ;
    END CO
    PIN CI
        AntennaGateArea              0.3780 ;
        AntennaPartialMetalArea      2.0434 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8108 LAYER met1 ;
    END CI
    PIN B
        AntennaGateArea              0.1260 ;
        AntennaPartialMetalArea      0.8553 LAYER met1 ;
        AntennaPartialMetalSideArea  0.7254 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.1260 ;
        AntennaPartialMetalArea      0.6058 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5238 LAYER met1 ;
    END A
    PIN GND
    END GND
END ADDFXL
MACRO ADDFX4
    PIN S
        AntennaPartialMetalArea      0.7960 LAYER met1 ;
        AntennaPartialMetalSideArea  0.4122 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END S
    PIN CO
        AntennaPartialMetalArea      1.2080 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5976 LAYER met1 ;
        AntennaDiffArea              1.4172 ;
    END CO
    PIN CI
        AntennaGateArea              0.3816 ;
        AntennaPartialMetalArea      1.9147 LAYER met1 ;
        AntennaPartialMetalSideArea  1.6776 LAYER met1 ;
    END CI
    PIN B
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.6492 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5382 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      1.2298 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8946 LAYER met1 ;
    END A
    PIN GND
    END GND
END ADDFX4
MACRO ADDFX2
    PIN S
        AntennaPartialMetalArea      1.1324 LAYER met1 ;
        AntennaPartialMetalSideArea  0.6966 LAYER met1 ;
        AntennaDiffArea              1.5600 ;
    END S
    PIN CO
        AntennaPartialMetalArea      0.8820 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5940 LAYER met1 ;
        AntennaDiffArea              1.5408 ;
    END CO
    PIN CI
        AntennaGateArea              0.3816 ;
        AntennaPartialMetalArea      2.0073 LAYER met1 ;
        AntennaPartialMetalSideArea  1.8000 LAYER met1 ;
    END CI
    PIN B
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.6492 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5382 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      1.2260 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8964 LAYER met1 ;
    END A
    PIN GND
    END GND
END ADDFX2
MACRO ADDFX1
    PIN S
        AntennaPartialMetalArea      0.7466 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5598 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END S
    PIN CO
        AntennaPartialMetalArea      0.7228 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5058 LAYER met1 ;
        AntennaDiffArea              0.7800 ;
    END CO
    PIN CI
        AntennaGateArea              0.3816 ;
        AntennaPartialMetalArea      2.0598 LAYER met1 ;
        AntennaPartialMetalSideArea  1.7550 LAYER met1 ;
    END CI
    PIN B
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      0.6512 LAYER met1 ;
        AntennaPartialMetalSideArea  0.5382 LAYER met1 ;
    END B
    PIN A
        AntennaGateArea              0.5400 ;
        AntennaPartialMetalArea      1.2260 LAYER met1 ;
        AntennaPartialMetalSideArea  0.8964 LAYER met1 ;
    END A
    PIN GND
    END GND
END ADDFX1
END LIBRARY
