#******
# Preview export LEF
#
#        Preview sub-version 4.4.2.100.41
#
# RC values have been extracted from UMC's worst case interconnect
# tables and worst case resistance values.
#
# Resistance and Capacitance Values
# ---------------------------------
# The LEF technology files included in this directory contain
# resistance and capacitance (RC) values for the purpose of timing
# driven place & route.  Please note that the RC values contained in
# this tech file were created using the worst case interconnect models
# from the foundry and assume a full metal route at every grid location
# on every metal layer, so the values are intentionally very
# conservative. It is assumed that this technology file will be used
# only as a starting point for creating initial timing driven place &
# route runs during the development of your own more accurate RC
# values, tailored to your specific place & route environment. AS A
# RESULT, TIMING NUMBERS DERIVED FROM THESE RC VALUES MAY BE
# SIGNIFICANTLY SLOWER THAN REALITY.
#
# The RC values used in the LEF technology file are to be used only
# for timing driven place & route. Due to accuracy limitations,
# please do not attempt to use this file for chip-level RC extraction
# in conjunction with your sign-off timing simulations. For chip-level
# extraction, please use a dedicated extraction tool such as HyperExtract,
# starRC or Simplex, etc.
#
# TECH LIB NAME: umc18
# TECH FILE NAME: techfile.cds
#
# $Id: umc18_6lm.lef,v 1.9 2003-11-18 17:09:25-08 prakash Exp $
#
#******    

VERSION 5.6 ;

NAMESCASESENSITIVE ON ;

UNITS
    DATABASE MICRONS 1000  ;
END UNITS

MANUFACTURINGGRID 0.01 ;

LAYER poly
    TYPE MASTERSLICE ;
END poly

LAYER met1
    TYPE ROUTING ;
    WIDTH 0.240 ;
    MAXWIDTH 9.0 ;
    AREA 0.1764 ;
    THICKNESS 0.528 ;
    SPACING 0.240 ;
    SPACING 0.240 RANGE 0.240 9.990 ;
    SPACING 0.280 RANGE 10.0 100000.0 ;
    PITCH 0.560 ;
    DIRECTION HORIZONTAL ;
    RESISTANCE RPERSQ 0.11500000 ;
    CAPACITANCE CPERSQDIST 1.3207e-04 ;
    EDGECAPACITANCE        8.7698e-05 ;
    ACCURRENTDENSITY AVERAGE 0.87 ;
    DCCURRENTDENSITY AVERAGE 0.87 ; 
END met1

LAYER via1
    TYPE CUT ;
    ACCURRENTDENSITY PEAK 67.0 ;
    DCCURRENTDENSITY AVERAGE 67.0 ;
END via1

LAYER met2
    TYPE ROUTING ;
    WIDTH 0.280 ;
    MAXWIDTH 9.0 ;
    AREA 0.1936 ;
    THICKNESS 0.638 ;
    SPACING 0.280 ;
    SPACING 0.280 RANGE 0.280 9.990 ;
    SPACING 0.320 RANGE 10.0 100000.0 ;
    PITCH 0.660 ;
    DIRECTION VERTICAL ;
    RESISTANCE RPERSQ 0.09500000 ;
    CAPACITANCE CPERSQDIST 7.0017e-05 ;
    EDGECAPACITANCE        8.3089e-05 ;
    ACCURRENTDENSITY AVERAGE 1.03 ;
    DCCURRENTDENSITY AVERAGE 1.03 ; 
END met2

LAYER via2
    TYPE CUT ;
    ACCURRENTDENSITY PEAK 67.0 ;
    DCCURRENTDENSITY AVERAGE 67.0 ;
END via2

LAYER met3
    TYPE ROUTING ;
    WIDTH 0.280 ;
    MAXWIDTH 9.0 ;
    AREA 0.1936 ;
    THICKNESS 0.638 ;
    SPACING 0.280 ;
    SPACING 0.280 RANGE 0.280 9.990 ;
    SPACING 0.320 RANGE 10.0 100000.0 ;
    PITCH 0.560 ;
    DIRECTION HORIZONTAL ;
    RESISTANCE RPERSQ 0.09500000 ;
    CAPACITANCE CPERSQDIST 6.3072e-05 ;
    EDGECAPACITANCE        1.0032e-04 ;
    ACCURRENTDENSITY AVERAGE 1.03 ;
    DCCURRENTDENSITY AVERAGE 1.03 ; 
END met3

LAYER via3
    TYPE CUT ;
    ACCURRENTDENSITY PEAK 67.0 ;
    DCCURRENTDENSITY AVERAGE 67.0 ;
END via3

LAYER met4
    TYPE ROUTING ;
    WIDTH 0.280 ;
    MAXWIDTH 9.0 ;
    AREA 0.1936 ; 
    THICKNESS 0.638 ;
    SPACING 0.280 ;
    SPACING 0.280 RANGE 0.280 9.990 ; 
    SPACING 0.320 RANGE 10.0 100000.0 ;
    PITCH 0.660 ;
    DIRECTION VERTICAL ;
    RESISTANCE RPERSQ 0.09500000 ;
    CAPACITANCE CPERSQDIST 5.9899e-05 ;
    EDGECAPACITANCE        8.2123e-05 ;
    ACCURRENTDENSITY AVERAGE 1.03 ;
    DCCURRENTDENSITY AVERAGE 1.03 ; 
END met4

LAYER via4
    TYPE CUT ;
    ACCURRENTDENSITY PEAK 67.0 ;
    DCCURRENTDENSITY AVERAGE 67.0 ;
END via4

LAYER met5
    TYPE ROUTING ;
    WIDTH 0.280 ;
    MAXWIDTH 9.0 ;
    AREA 0.1936 ;
    THICKNESS 0.6380 ;
    SPACING 0.280 ;
    SPACING 0.280 RANGE 0.280 9.990 ;
    SPACING 0.320 RANGE 10.0 100000.0 ;
    PITCH 0.560 ;
    DIRECTION HORIZONTAL ;
    RESISTANCE RPERSQ 0.09500000 ;
    CAPACITANCE CPERSQDIST 4.8187e-05 ;
    EDGECAPACITANCE        5.7617e-05 ;
    ACCURRENTDENSITY AVERAGE 1.03 ;
    DCCURRENTDENSITY AVERAGE 1.03 ; 
END met5

LAYER via5
    TYPE CUT ;
    ACCURRENTDENSITY PEAK 67.0 ;
    DCCURRENTDENSITY AVERAGE 67.0 ;
END via5

LAYER met6
    TYPE ROUTING ;
    WIDTH 0.440 ;
    MAXWIDTH 9.0 ;
    AREA 0.4624 ;
    THICKNESS 0.9460 ;
    SPACING 0.440 ;
    SPACING 0.440 RANGE 0.440 9.990 ;
    SPACING 0.600 RANGE 10.0 100000.0 ;
    PITCH 1.320 ;
    DIRECTION VERTICAL ;
    RESISTANCE RPERSQ 0.05500000 ;
    CAPACITANCE CPERSQDIST 2.5901e-05 ;
    EDGECAPACITANCE        8.5684e-05 ;
    ACCURRENTDENSITY AVERAGE 1.74 ;
    DCCURRENTDENSITY AVERAGE 1.74 ; 
END met6

LAYER OVERLAP
    TYPE OVERLAP ;
END OVERLAP

VIA Via1 DEFAULT
    # Worst case via resistance
    RESISTANCE 15.000e+00 ;
    LAYER met1 ;
        RECT -0.220 -0.140 0.220 0.140 ;
    LAYER via1 ;
        RECT -0.140 -0.140 0.140 0.140 ;
    LAYER met2 ;
        RECT -0.220 -0.140 0.220 0.140 ;
END Via1

VIA Via2 DEFAULT
    # Worst case via resistance
    RESISTANCE 15.000e+00 ;
    LAYER met2 ;
        RECT -0.220 -0.140 0.220 0.140 ;
    LAYER via2 ;
        RECT -0.140 -0.140 0.140 0.140 ;
    LAYER met3 ;
        RECT -0.220 -0.140 0.220 0.140 ;
END Via2

VIA Via2ts DEFAULT TOPOFSTACKONLY
    # Worst case via resistance
    RESISTANCE 15.000e+00 ;
    LAYER met2 ;
        RECT -0.220 -0.140 0.220 0.300 ;
    LAYER via2 ;
        RECT -0.140 -0.140 0.140 0.140 ;
    LAYER met3 ;
        RECT -0.220 -0.140 0.220 0.140 ;
END Via2ts

VIA Via3 DEFAULT
    # Worst case via resistance
    RESISTANCE 15.000e+00 ;
    LAYER met3 ;
        RECT -0.220 -0.140 0.220 0.140 ;
    LAYER via3 ;
        RECT -0.140 -0.140 0.140 0.140 ;
    LAYER met4 ;
        RECT -0.220 -0.140 0.220 0.140 ;
END Via3

VIA Via3ts DEFAULT TOPOFSTACKONLY
    # Worst case via resistance
    RESISTANCE 15.000e+00 ;
    LAYER met3 ;
        RECT -0.220 -0.140 0.220 0.300 ;
    LAYER via3 ;
        RECT -0.140 -0.140 0.140 0.140 ;
    LAYER met4 ;
        RECT -0.220 -0.140 0.220 0.140 ;
END Via3ts

VIA Via4 DEFAULT
    # Worst case via resistance
    RESISTANCE 15.000e+00 ;
    LAYER met4 ;
        RECT -0.220 -0.140 0.220 0.140 ;
    LAYER via4 ;
        RECT -0.140 -0.140 0.140 0.140 ;
    LAYER met5 ;
        RECT -0.220 -0.140 0.220 0.140 ;
END Via4

VIA Via4ts DEFAULT TOPOFSTACKONLY
    # Worst case via resistance
    RESISTANCE 15.000e+00 ;
    LAYER met4 ;
        RECT -0.220 -0.140 0.220 0.300 ;
    LAYER via4 ;
        RECT -0.140 -0.140 0.140 0.140 ;
    LAYER met5 ;
        RECT -0.220 -0.140 0.220 0.140 ;
END Via4ts

VIA Via5 DEFAULT
    # Worst case via resistance
    RESISTANCE 15.000e+00 ;
    LAYER met5 ;
        RECT -0.220 -0.140 0.220 0.140 ;
    LAYER via5 ;
        RECT -0.140 -0.140 0.140 0.140 ;
    LAYER met6 ;
        RECT -0.260 -0.220 0.260 0.220 ;
END Via5

VIA Via5ts DEFAULT TOPOFSTACKONLY
    # Worst case via resistance
    RESISTANCE 15.000e+00 ;
    LAYER met5 ;
        RECT -0.220 -0.140 0.220 0.300 ;
    LAYER via5 ;
        RECT -0.140 -0.140 0.140 0.140 ;
    LAYER met6 ;
        RECT -0.260 -0.220 0.260 0.220 ;
END Via5ts

VIARULE via1Array GENERATE
    LAYER met1 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.20 ;
        METALOVERHANG 0.000 ;

    LAYER met2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.20 ;
        METALOVERHANG 0.000 ;

    LAYER via1 ;
        RECT -0.140 -0.140 0.140 0.140 ;
        SPACING 0.560 BY 0.560 ;
END via1Array

VIARULE via2Array GENERATE
    LAYER met2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.20 ;
        METALOVERHANG 0.000 ;

    LAYER met3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.20 ;
        METALOVERHANG 0.000 ;

    LAYER via2 ;
        RECT -0.140 -0.140 0.140 0.140 ;
        SPACING 0.560 BY 0.560 ;
END via2Array

VIARULE via3Array GENERATE
    LAYER met3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.20 ;
        METALOVERHANG 0.000 ;

    LAYER met4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.20 ;
        METALOVERHANG 0.000 ;

    LAYER via3 ;
        RECT -0.140 -0.140 0.140 0.140 ;
        SPACING 0.560 BY 0.560 ;
END via3Array

VIARULE via4Array GENERATE
    LAYER met4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.20 ;
        METALOVERHANG 0.000 ;

    LAYER met5 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.20 ;
        METALOVERHANG 0.000 ;

    LAYER via4 ;
        RECT -0.140 -0.140 0.140 0.140 ;
        SPACING 0.560 BY 0.560 ;
END via4Array

VIARULE via5Array GENERATE
    LAYER met5 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.20 ;
        METALOVERHANG 0.000 ;

    LAYER met6 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.20 ;
        METALOVERHANG 0.000 ;

    LAYER via5 ;
        RECT -0.140 -0.140 0.140 0.140 ;
        SPACING 0.560 BY 0.560 ;
END via5Array

VIARULE TURNM1 GENERATE
    LAYER met1 ;
        DIRECTION vertical ;

    LAYER met1 ;
        DIRECTION horizontal ;
END TURNM1

VIARULE TURNM2 GENERATE
    LAYER met2 ;
        DIRECTION vertical ;

    LAYER met2 ;
        DIRECTION horizontal ;
END TURNM2

VIARULE TURNM3 GENERATE
    LAYER met3 ;
        DIRECTION vertical ;

    LAYER met3 ;
        DIRECTION horizontal ;
END TURNM3

VIARULE TURNM4 GENERATE
    LAYER met4 ;
        DIRECTION vertical ;

    LAYER met4 ;
        DIRECTION horizontal ;
END TURNM4

VIARULE TURNM5 GENERATE
    LAYER met5 ;
        DIRECTION vertical ;

    LAYER met5 ;
        DIRECTION horizontal ;
END TURNM5

VIARULE TURNM6 GENERATE
    LAYER met6 ;
        DIRECTION vertical ;

    LAYER met6 ;
        DIRECTION horizontal ;
END TURNM6

SPACING
    SAMENET met1 met1 0.240  ;
    SAMENET met2 met2 0.280  STACK ;
    SAMENET met3 met3 0.280  STACK ;
    SAMENET met4 met4 0.280  STACK ;
    SAMENET met5 met5 0.280  STACK ;
    SAMENET met6 met6 0.440  STACK ;
    SAMENET via1 via1 0.280  ;
    SAMENET via2 via2 0.280  ;
    SAMENET via3 via3 0.280  ;
    SAMENET via4 via4 0.280  ;
    SAMENET via5 via5 0.280  ;
    SAMENET via1 via2 0.000  STACK ;
    SAMENET via2 via3 0.000  STACK ;
    SAMENET via3 via4 0.000  STACK ;
    SAMENET via4 via5 0.000  STACK ;
END SPACING

SITE umc6site
    SYMMETRY y  ;
    CLASS CORE ;
    SIZE 0.660 BY 5.040 ;
END umc6site

MACRO RFRDX4
    CLASS CORE ;
    FOREIGN RFRDX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.460 2.060 1.860 2.460 ;
        RECT  1.860 2.060 2.830 2.300 ;
        RECT  2.830 1.580 2.850 2.300 ;
        RECT  2.850 1.580 2.900 2.400 ;
        RECT  2.900 1.580 3.090 3.480 ;
        RECT  3.090 1.420 3.300 3.480 ;
        RECT  3.300 1.420 3.800 1.820 ;
        END
    END RB
    PIN BRB
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.770 1.820 0.880 3.220 ;
        RECT  0.880 0.920 1.210 4.120 ;
        RECT  1.210 2.700 1.280 4.120 ;
        RECT  1.210 0.920 1.280 1.820 ;
        RECT  1.280 2.700 1.530 3.220 ;
        RECT  1.530 2.700 2.210 2.960 ;
        RECT  2.210 2.540 2.610 2.960 ;
        END
    END BRB
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.080 0.530 5.440 ;
        RECT  0.530 3.780 0.560 5.440 ;
        RECT  0.560 4.640 1.600 5.440 ;
        RECT  1.600 3.580 2.000 5.440 ;
        RECT  2.000 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 1.560 ;
        RECT  0.560 -0.400 1.600 0.400 ;
        RECT  1.600 -0.400 2.000 1.060 ;
        RECT  2.000 -0.400 3.960 0.400 ;
        END
    END GND
END RFRDX4

MACRO RFRDX2
    CLASS CORE ;
    FOREIGN RFRDX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ RFRDX4 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.650 2.060 1.050 2.460 ;
        RECT  1.050 2.060 2.170 2.300 ;
        RECT  2.170 1.580 2.180 2.300 ;
        RECT  2.180 1.580 2.430 3.480 ;
        RECT  2.430 1.420 2.580 3.480 ;
        RECT  2.580 1.420 3.140 1.820 ;
        END
    END RB
    PIN BRB
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.160 0.920 0.400 4.120 ;
        RECT  0.400 2.720 0.560 4.120 ;
        RECT  0.400 0.920 0.560 1.820 ;
        RECT  0.560 2.940 1.490 3.220 ;
        RECT  1.490 2.540 1.750 3.220 ;
        RECT  1.750 2.540 1.890 2.960 ;
        END
    END BRB
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.880 5.440 ;
        RECT  0.880 3.580 1.280 5.440 ;
        RECT  1.280 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.880 0.400 ;
        RECT  0.880 -0.400 1.280 1.560 ;
        RECT  1.280 -0.400 3.300 0.400 ;
        END
    END GND
END RFRDX2

MACRO RFRDX1
    CLASS CORE ;
    FOREIGN RFRDX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ RFRDX4 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.650 2.060 1.050 2.460 ;
        RECT  1.050 2.060 2.170 2.300 ;
        RECT  2.170 1.580 2.180 2.300 ;
        RECT  2.180 1.580 2.430 3.480 ;
        RECT  2.430 1.420 2.580 3.480 ;
        RECT  2.580 1.420 3.140 1.820 ;
        END
    END RB
    PIN BRB
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.160 1.420 0.400 3.480 ;
        RECT  0.400 2.940 0.560 3.480 ;
        RECT  0.400 1.420 0.560 1.820 ;
        RECT  0.560 2.940 1.490 3.220 ;
        RECT  1.490 2.540 1.750 3.220 ;
        RECT  1.750 2.540 1.890 2.960 ;
        END
    END BRB
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.880 5.440 ;
        RECT  0.880 3.540 1.280 5.440 ;
        RECT  1.280 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.880 0.400 ;
        RECT  0.880 -0.400 1.280 1.740 ;
        RECT  1.280 -0.400 3.300 0.400 ;
        END
    END GND
END RFRDX1

MACRO RF2R1WX2
    CLASS CORE ;
    FOREIGN RF2R1WX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN WW
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.710 2.060 0.950 2.460 ;
        RECT  0.950 2.140 1.520 2.380 ;
        RECT  1.520 2.140 1.760 3.710 ;
        RECT  1.760 2.140 1.800 2.400 ;
        RECT  1.800 1.890 1.870 2.400 ;
        RECT  1.760 3.470 2.120 3.710 ;
        RECT  1.870 1.890 2.200 2.380 ;
        RECT  2.120 3.470 2.300 3.780 ;
        RECT  2.300 3.470 2.540 4.140 ;
        RECT  2.540 3.740 2.700 4.140 ;
        END
    END WW
    PIN WB
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.460 0.660 1.780 1.530 ;
        RECT  1.780 0.660 1.860 0.900 ;
        END
    END WB
    PIN R2W
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.460 1.830 7.520 2.090 ;
        RECT  7.520 1.830 7.720 2.480 ;
        RECT  7.720 1.840 7.810 2.480 ;
        RECT  7.810 2.080 7.920 2.480 ;
        END
    END R2W
    PIN R2B
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  8.750 2.820 8.920 3.720 ;
        RECT  8.780 0.920 8.920 1.820 ;
        RECT  8.920 0.920 9.160 3.720 ;
        RECT  9.160 0.920 9.180 1.820 ;
        END
    END R2B
    PIN R1W
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.460 0.640 7.120 1.040 ;
        END
    END R1W
    PIN R1B
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  5.480 1.270 5.730 1.530 ;
        RECT  5.730 0.920 5.760 1.530 ;
        RECT  5.760 0.920 6.000 3.620 ;
        RECT  6.000 2.720 6.160 3.620 ;
        RECT  6.000 0.920 6.220 1.820 ;
        END
    END R1B
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.750 5.440 ;
        RECT  0.750 4.430 1.150 5.440 ;
        RECT  1.150 4.640 3.320 5.440 ;
        RECT  3.320 4.480 3.720 5.440 ;
        RECT  3.720 4.640 4.510 5.440 ;
        RECT  4.510 3.900 4.940 5.440 ;
        RECT  4.940 4.640 7.270 5.440 ;
        RECT  7.270 3.900 7.670 5.440 ;
        RECT  7.670 4.640 10.000 5.440 ;
        RECT  10.000 2.890 10.400 5.440 ;
        RECT  10.400 4.640 10.560 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.820 0.400 ;
        RECT  0.820 -0.400 1.220 0.610 ;
        RECT  1.220 -0.400 3.260 0.400 ;
        RECT  3.260 -0.400 3.660 1.100 ;
        RECT  3.660 -0.400 4.570 0.400 ;
        RECT  4.570 -0.400 4.970 0.610 ;
        RECT  4.970 -0.400 7.400 0.400 ;
        RECT  7.400 -0.400 7.800 0.610 ;
        RECT  7.800 -0.400 10.000 0.400 ;
        RECT  10.000 -0.400 10.400 1.560 ;
        RECT  10.400 -0.400 10.560 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  9.750 2.070 10.120 2.470 ;
        RECT  9.720 2.070 9.750 4.210 ;
        RECT  9.510 2.230 9.720 4.210 ;
        RECT  8.290 3.970 9.510 4.210 ;
        RECT  8.500 2.180 8.680 2.580 ;
        RECT  8.400 1.420 8.500 2.580 ;
        RECT  8.160 1.420 8.400 3.120 ;
        RECT  8.050 3.420 8.290 4.210 ;
        RECT  8.060 1.420 8.160 1.820 ;
        RECT  7.970 2.720 8.160 3.120 ;
        RECT  6.650 3.420 8.050 3.660 ;
        RECT  6.720 1.420 6.940 1.820 ;
        RECT  6.720 2.720 6.880 3.120 ;
        RECT  6.540 1.420 6.720 3.120 ;
        RECT  6.410 3.420 6.650 4.100 ;
        RECT  6.480 1.500 6.540 3.120 ;
        RECT  6.240 2.060 6.480 2.460 ;
        RECT  5.520 3.860 6.410 4.100 ;
        RECT  5.280 2.440 5.520 4.100 ;
        RECT  5.180 2.440 5.280 2.680 ;
        RECT  4.680 2.180 5.180 2.680 ;
        RECT  4.450 1.380 4.680 2.680 ;
        RECT  4.440 1.300 4.450 2.680 ;
        RECT  4.050 1.300 4.440 1.700 ;
        RECT  4.430 2.440 4.440 2.680 ;
        RECT  4.030 2.440 4.430 3.300 ;
        RECT  2.680 1.940 4.200 2.180 ;
        RECT  3.120 2.440 4.030 2.680 ;
        RECT  2.540 1.330 2.680 3.200 ;
        RECT  2.440 1.250 2.540 3.200 ;
        RECT  2.140 1.250 2.440 1.650 ;
        RECT  2.000 2.960 2.440 3.200 ;
        RECT  1.450 3.950 1.850 4.350 ;
        RECT  0.560 3.950 1.450 4.190 ;
        RECT  0.400 1.320 0.560 1.720 ;
        RECT  0.400 2.720 0.560 4.190 ;
        RECT  0.320 1.320 0.400 4.190 ;
        RECT  0.160 1.320 0.320 3.120 ;
    END
END RF2R1WX2

MACRO RF1R1WX2
    CLASS CORE ;
    FOREIGN RF1R1WX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN WW
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.360 0.920 2.760 ;
        RECT  0.920 2.360 1.460 2.600 ;
        RECT  1.460 2.360 1.530 2.660 ;
        RECT  1.530 2.360 1.770 3.700 ;
        RECT  1.770 2.360 1.810 2.660 ;
        RECT  1.810 1.580 2.050 2.660 ;
        RECT  2.050 1.580 2.210 1.980 ;
        RECT  1.770 3.460 2.330 3.700 ;
        RECT  2.330 3.460 2.730 3.860 ;
        END
    END WW
    PIN WB
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 1.090 2.090 ;
        RECT  1.090 1.680 1.120 2.090 ;
        RECT  1.120 1.680 1.490 2.080 ;
        END
    END WB
    PIN RWN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.400 4.000 4.830 4.400 ;
        RECT  4.830 4.000 6.050 4.240 ;
        RECT  6.050 3.500 6.290 4.240 ;
        RECT  6.290 3.500 6.460 3.780 ;
        END
    END RWN
    PIN RW
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.870 0.640 4.350 1.010 ;
        RECT  4.350 0.640 4.590 1.040 ;
        END
    END RW
    PIN RB
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  4.730 2.640 4.890 3.120 ;
        RECT  4.820 1.830 4.890 2.090 ;
        RECT  4.890 0.780 5.130 3.120 ;
        END
    END RB
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.750 5.440 ;
        RECT  0.750 4.420 1.150 5.440 ;
        RECT  1.150 4.640 3.180 5.440 ;
        RECT  3.180 3.520 3.580 5.440 ;
        RECT  3.580 4.640 6.040 5.440 ;
        RECT  6.040 4.480 6.440 5.440 ;
        RECT  6.440 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.030 0.400 ;
        RECT  1.030 -0.400 1.430 0.630 ;
        RECT  1.430 -0.400 3.220 0.400 ;
        RECT  3.220 -0.400 3.620 1.060 ;
        RECT  3.620 -0.400 5.990 0.400 ;
        RECT  5.990 -0.400 6.390 1.420 ;
        RECT  6.390 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.650 1.900 6.140 2.140 ;
        RECT  5.410 1.900 5.650 3.600 ;
        RECT  4.480 3.360 5.410 3.600 ;
        RECT  4.240 1.300 4.480 3.600 ;
        RECT  4.080 1.300 4.240 1.700 ;
        RECT  3.970 2.900 4.240 3.300 ;
        RECT  3.800 1.940 4.000 2.340 ;
        RECT  3.320 2.900 3.970 3.140 ;
        RECT  3.560 1.880 3.800 2.340 ;
        RECT  2.690 1.880 3.560 2.120 ;
        RECT  3.080 2.360 3.320 3.140 ;
        RECT  2.450 0.940 2.690 3.220 ;
        RECT  2.170 0.940 2.450 1.340 ;
        RECT  2.020 2.980 2.450 3.220 ;
        RECT  1.510 3.940 1.910 4.400 ;
        RECT  0.560 3.940 1.510 4.180 ;
        RECT  0.400 0.720 0.560 1.120 ;
        RECT  0.400 3.000 0.560 4.180 ;
        RECT  0.320 0.720 0.400 4.180 ;
        RECT  0.160 0.720 0.320 3.400 ;
    END
END RF1R1WX2

MACRO AFCSHCONX4
    CLASS CORE ;
    FOREIGN AFCSHCONX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 38.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  38.410 1.520 38.510 3.150 ;
        RECT  38.290 0.870 38.410 3.150 ;
        RECT  38.270 0.870 38.290 4.250 ;
        RECT  38.170 0.870 38.270 2.100 ;
        RECT  38.050 2.850 38.270 4.250 ;
        RECT  37.730 0.700 38.170 2.100 ;
        END
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  36.450 1.820 36.850 2.400 ;
        RECT  36.410 1.820 36.450 2.100 ;
        END
    END CS
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  22.550 2.210 25.800 2.450 ;
        RECT  22.650 3.650 25.670 3.890 ;
        RECT  22.330 3.500 22.650 3.890 ;
        RECT  22.330 2.210 22.550 2.760 ;
        RECT  21.890 2.210 22.330 3.890 ;
        END
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.260 2.240 21.420 4.400 ;
        RECT  21.180 1.600 21.260 4.400 ;
        RECT  21.020 1.600 21.180 2.480 ;
        RECT  19.340 4.160 21.180 4.400 ;
        RECT  20.790 1.600 21.020 1.840 ;
        RECT  19.110 3.720 19.340 4.400 ;
        RECT  19.100 3.190 19.110 4.400 ;
        RECT  19.030 3.190 19.100 3.990 ;
        RECT  18.870 2.380 19.030 3.990 ;
        RECT  18.830 2.380 18.870 3.780 ;
        RECT  18.590 2.080 18.830 3.780 ;
        RECT  18.430 2.080 18.590 3.430 ;
        RECT  17.760 3.190 18.430 3.430 ;
        RECT  17.520 3.190 17.760 3.700 ;
        END
    END CO0N
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  30.760 2.340 31.660 2.740 ;
        END
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  11.090 2.370 12.490 2.770 ;
        END
    END CI0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.560 2.250 5.960 2.740 ;
        RECT  5.470 2.260 5.560 2.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.190 2.380 1.210 3.220 ;
        RECT  0.790 2.120 1.190 3.220 ;
        RECT  0.770 2.380 0.790 3.220 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  37.600 4.640 38.940 5.440 ;
        RECT  37.200 3.910 37.600 5.440 ;
        RECT  36.660 4.640 37.200 5.440 ;
        RECT  36.420 3.860 36.660 5.440 ;
        RECT  32.980 4.640 36.420 5.440 ;
        RECT  32.580 3.320 32.980 5.440 ;
        RECT  31.540 4.640 32.580 5.440 ;
        RECT  31.140 4.080 31.540 5.440 ;
        RECT  30.020 4.640 31.140 5.440 ;
        RECT  29.780 4.080 30.020 5.440 ;
        RECT  13.770 4.640 29.780 5.440 ;
        RECT  13.370 4.480 13.770 5.440 ;
        RECT  12.150 4.640 13.370 5.440 ;
        RECT  11.750 4.480 12.150 5.440 ;
        RECT  10.850 4.640 11.750 5.440 ;
        RECT  10.450 4.480 10.850 5.440 ;
        RECT  9.270 4.640 10.450 5.440 ;
        RECT  8.870 4.480 9.270 5.440 ;
        RECT  6.350 4.640 8.870 5.440 ;
        RECT  5.950 4.480 6.350 5.440 ;
        RECT  2.510 4.640 5.950 5.440 ;
        RECT  2.110 4.080 2.510 5.440 ;
        RECT  1.280 4.640 2.110 5.440 ;
        RECT  0.880 4.060 1.280 5.440 ;
        RECT  0.000 4.640 0.880 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  37.490 -0.400 38.940 0.400 ;
        RECT  37.090 -0.400 37.490 0.610 ;
        RECT  36.020 -0.400 37.090 0.400 ;
        RECT  35.780 -0.400 36.020 1.820 ;
        RECT  32.910 -0.400 35.780 0.400 ;
        RECT  32.510 -0.400 32.910 0.560 ;
        RECT  31.330 -0.400 32.510 0.400 ;
        RECT  30.930 -0.400 31.330 0.560 ;
        RECT  29.740 -0.400 30.930 0.400 ;
        RECT  29.340 -0.400 29.740 0.560 ;
        RECT  14.130 -0.400 29.340 0.400 ;
        RECT  13.730 -0.400 14.130 0.980 ;
        RECT  9.690 -0.400 13.730 0.400 ;
        RECT  9.290 -0.400 9.690 0.840 ;
        RECT  8.110 -0.400 9.290 0.400 ;
        RECT  7.710 -0.400 8.110 0.560 ;
        RECT  2.630 -0.400 7.710 0.400 ;
        RECT  2.230 -0.400 2.630 0.560 ;
        RECT  1.280 -0.400 2.230 0.400 ;
        RECT  0.880 -0.400 1.280 1.560 ;
        RECT  0.000 -0.400 0.880 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  37.810 2.340 37.970 2.580 ;
        RECT  37.570 2.340 37.810 3.600 ;
        RECT  36.180 3.360 37.570 3.600 ;
        RECT  37.090 1.340 37.330 3.120 ;
        RECT  36.520 1.340 37.090 1.580 ;
        RECT  35.700 2.880 37.090 3.120 ;
        RECT  35.940 3.360 36.180 4.370 ;
        RECT  34.100 4.130 35.940 4.370 ;
        RECT  35.540 2.060 35.700 2.460 ;
        RECT  35.460 2.880 35.700 3.890 ;
        RECT  35.300 0.800 35.540 2.460 ;
        RECT  34.580 3.650 35.460 3.890 ;
        RECT  26.740 0.800 35.300 1.040 ;
        RECT  35.060 3.170 35.220 3.410 ;
        RECT  34.820 1.370 35.060 3.410 ;
        RECT  34.340 2.140 34.580 3.890 ;
        RECT  34.100 1.350 34.420 1.750 ;
        RECT  33.860 1.350 34.100 4.370 ;
        RECT  33.380 1.330 33.620 4.220 ;
        RECT  32.900 1.280 33.140 2.700 ;
        RECT  28.160 1.280 32.900 1.520 ;
        RECT  32.180 3.300 32.260 4.200 ;
        RECT  31.940 1.760 32.180 4.200 ;
        RECT  31.720 1.760 31.940 2.000 ;
        RECT  31.860 3.300 31.940 4.200 ;
        RECT  29.540 3.600 31.860 3.840 ;
        RECT  30.450 3.100 30.820 3.340 ;
        RECT  30.450 1.760 30.530 2.000 ;
        RECT  30.130 1.760 30.450 3.340 ;
        RECT  29.290 3.100 30.130 3.340 ;
        RECT  29.300 3.600 29.540 4.400 ;
        RECT  26.440 4.160 29.300 4.400 ;
        RECT  29.060 2.350 29.290 3.340 ;
        RECT  29.050 2.350 29.060 3.920 ;
        RECT  28.820 3.100 29.050 3.920 ;
        RECT  28.720 1.760 28.950 2.000 ;
        RECT  27.220 3.680 28.820 3.920 ;
        RECT  28.580 1.760 28.720 2.810 ;
        RECT  28.480 1.760 28.580 3.440 ;
        RECT  28.340 2.570 28.480 3.440 ;
        RECT  28.180 3.200 28.340 3.440 ;
        RECT  28.000 1.280 28.160 1.840 ;
        RECT  27.870 1.280 28.000 2.910 ;
        RECT  27.760 1.280 27.870 3.440 ;
        RECT  27.630 2.670 27.760 3.440 ;
        RECT  27.460 3.200 27.630 3.440 ;
        RECT  27.220 1.440 27.440 1.840 ;
        RECT  26.980 1.440 27.220 3.920 ;
        RECT  26.700 3.440 26.980 3.840 ;
        RECT  26.500 0.800 26.740 1.970 ;
        RECT  21.740 1.730 26.500 1.970 ;
        RECT  26.200 2.930 26.440 4.400 ;
        RECT  26.020 0.740 26.260 1.140 ;
        RECT  22.780 2.930 26.200 3.170 ;
        RECT  22.460 0.740 26.020 0.980 ;
        RECT  22.220 1.250 25.580 1.490 ;
        RECT  21.980 0.640 22.220 1.490 ;
        RECT  14.610 0.640 21.980 0.880 ;
        RECT  21.500 1.120 21.740 1.970 ;
        RECT  20.550 1.120 21.500 1.360 ;
        RECT  20.780 2.720 20.940 3.920 ;
        RECT  20.700 2.280 20.780 3.920 ;
        RECT  20.550 2.280 20.700 2.960 ;
        RECT  19.820 3.680 20.700 3.920 ;
        RECT  20.540 1.120 20.550 2.960 ;
        RECT  20.310 1.120 20.540 2.520 ;
        RECT  20.300 3.200 20.460 3.440 ;
        RECT  20.070 2.760 20.300 3.440 ;
        RECT  20.060 2.240 20.070 3.440 ;
        RECT  19.990 2.240 20.060 3.000 ;
        RECT  19.830 1.120 19.990 3.000 ;
        RECT  19.750 1.120 19.830 2.480 ;
        RECT  19.590 3.240 19.820 3.920 ;
        RECT  15.090 1.120 19.750 1.360 ;
        RECT  19.580 2.720 19.590 3.920 ;
        RECT  19.510 2.720 19.580 3.480 ;
        RECT  19.350 1.600 19.510 3.480 ;
        RECT  19.270 1.600 19.350 2.960 ;
        RECT  16.210 1.600 19.270 1.840 ;
        RECT  17.280 4.020 18.630 4.260 ;
        RECT  17.910 2.080 18.110 2.320 ;
        RECT  17.670 2.080 17.910 2.800 ;
        RECT  17.280 2.560 17.670 2.800 ;
        RECT  16.690 2.080 17.390 2.320 ;
        RECT  17.040 2.560 17.280 4.400 ;
        RECT  14.250 4.160 17.040 4.400 ;
        RECT  16.690 3.040 16.800 3.920 ;
        RECT  16.560 2.080 16.690 3.920 ;
        RECT  16.450 2.080 16.560 3.280 ;
        RECT  14.730 3.680 16.560 3.920 ;
        RECT  16.130 1.600 16.210 2.820 ;
        RECT  15.970 1.600 16.130 3.440 ;
        RECT  15.890 2.580 15.970 3.440 ;
        RECT  15.690 3.200 15.890 3.440 ;
        RECT  15.650 1.600 15.730 1.840 ;
        RECT  15.410 1.600 15.650 2.940 ;
        RECT  15.330 1.600 15.410 1.840 ;
        RECT  15.370 2.700 15.410 2.940 ;
        RECT  15.130 2.700 15.370 3.440 ;
        RECT  14.070 2.180 15.170 2.420 ;
        RECT  14.970 3.200 15.130 3.440 ;
        RECT  14.850 1.120 15.090 1.940 ;
        RECT  13.070 1.700 14.850 1.940 ;
        RECT  14.490 3.520 14.730 3.920 ;
        RECT  14.370 0.640 14.610 1.460 ;
        RECT  14.070 3.520 14.490 3.760 ;
        RECT  11.410 1.220 14.370 1.460 ;
        RECT  14.010 4.000 14.250 4.400 ;
        RECT  13.830 2.180 14.070 3.760 ;
        RECT  3.080 4.000 14.010 4.240 ;
        RECT  13.670 2.560 13.830 2.960 ;
        RECT  11.640 3.520 13.830 3.760 ;
        RECT  10.170 0.740 13.470 0.980 ;
        RECT  12.830 1.700 13.070 3.280 ;
        RECT  11.900 1.700 12.830 1.940 ;
        RECT  12.540 3.040 12.830 3.280 ;
        RECT  10.430 3.330 11.640 3.760 ;
        RECT  11.170 1.220 11.410 1.820 ;
        RECT  6.980 1.580 11.170 1.820 ;
        RECT  10.430 2.060 10.790 2.300 ;
        RECT  10.190 2.060 10.430 3.760 ;
        RECT  9.660 3.330 10.190 3.730 ;
        RECT  9.930 0.740 10.170 1.340 ;
        RECT  7.460 1.100 9.930 1.340 ;
        RECT  8.840 2.060 9.080 3.740 ;
        RECT  8.180 2.060 8.840 2.460 ;
        RECT  4.060 3.500 8.840 3.740 ;
        RECT  8.070 2.720 8.470 3.260 ;
        RECT  6.490 3.020 8.070 3.260 ;
        RECT  7.220 0.640 7.460 1.340 ;
        RECT  6.980 2.540 7.300 2.780 ;
        RECT  6.280 0.640 7.220 0.880 ;
        RECT  6.740 1.160 6.980 2.780 ;
        RECT  6.730 1.160 6.740 1.820 ;
        RECT  6.580 1.160 6.730 1.400 ;
        RECT  6.280 1.710 6.490 3.260 ;
        RECT  6.250 0.640 6.280 3.260 ;
        RECT  6.040 0.640 6.250 1.950 ;
        RECT  5.140 3.020 5.560 3.260 ;
        RECT  5.140 1.380 5.470 1.780 ;
        RECT  4.900 1.380 5.140 3.260 ;
        RECT  4.550 0.660 4.950 1.060 ;
        RECT  4.780 2.030 4.900 2.430 ;
        RECT  4.540 2.750 4.590 3.150 ;
        RECT  4.540 0.820 4.550 1.060 ;
        RECT  4.300 0.820 4.540 3.150 ;
        RECT  2.020 0.820 4.300 1.060 ;
        RECT  3.820 1.380 4.060 3.740 ;
        RECT  3.550 2.840 3.820 3.740 ;
        RECT  3.260 1.380 3.420 1.780 ;
        RECT  3.020 1.380 3.260 3.120 ;
        RECT  2.840 3.570 3.080 4.240 ;
        RECT  2.830 2.720 3.020 3.120 ;
        RECT  0.480 3.570 2.840 3.810 ;
        RECT  2.350 2.070 2.750 2.470 ;
        RECT  2.020 2.110 2.350 2.460 ;
        RECT  1.780 0.820 2.020 3.120 ;
        RECT  1.600 1.420 1.780 1.820 ;
        RECT  1.600 2.720 1.780 3.120 ;
        RECT  0.480 0.900 0.560 1.800 ;
        RECT  0.240 0.900 0.480 4.320 ;
        RECT  0.160 0.900 0.240 1.800 ;
    END
END AFCSHCONX4

MACRO AFCSHCONX2
    CLASS CORE ;
    FOREIGN AFCSHCONX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AFCSHCONX4 ;
    SIZE 35.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  35.240 0.840 35.480 4.370 ;
        RECT  35.080 0.840 35.240 1.740 ;
        RECT  35.080 2.970 35.240 4.370 ;
        RECT  34.430 1.260 35.080 1.540 ;
        END
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  33.150 1.820 33.550 2.360 ;
        END
    END CS
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  20.670 2.210 23.550 2.450 ;
        RECT  20.670 3.650 21.480 3.890 ;
        RECT  20.620 2.210 20.670 2.660 ;
        RECT  20.620 3.500 20.670 3.890 ;
        RECT  20.380 2.210 20.620 3.890 ;
        RECT  19.910 2.380 20.380 3.220 ;
        END
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  19.900 3.550 20.140 4.400 ;
        RECT  18.060 4.160 19.900 4.400 ;
        RECT  17.820 3.220 18.060 4.400 ;
        RECT  17.710 3.220 17.820 3.460 ;
        RECT  17.690 2.380 17.710 3.460 ;
        RECT  17.290 2.080 17.690 3.460 ;
        RECT  17.270 2.380 17.290 3.460 ;
        RECT  16.620 3.220 17.270 3.460 ;
        RECT  16.380 3.220 16.620 3.920 ;
        END
    END CO0N
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  28.580 2.390 28.840 2.700 ;
        RECT  27.840 2.460 28.580 2.700 ;
        END
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  11.110 2.370 11.370 2.770 ;
        RECT  10.790 2.370 11.110 3.220 ;
        RECT  10.760 2.950 10.790 3.210 ;
        END
    END CI0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.560 2.250 5.960 2.740 ;
        RECT  5.470 2.260 5.560 2.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.190 2.380 1.210 3.220 ;
        RECT  0.790 2.120 1.190 3.220 ;
        RECT  0.770 2.380 0.790 3.220 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  34.760 4.640 35.640 5.440 ;
        RECT  34.360 3.840 34.760 5.440 ;
        RECT  33.820 4.640 34.360 5.440 ;
        RECT  33.580 3.860 33.820 5.440 ;
        RECT  30.140 4.640 33.580 5.440 ;
        RECT  29.740 3.370 30.140 5.440 ;
        RECT  27.770 4.640 29.740 5.440 ;
        RECT  27.530 4.140 27.770 5.440 ;
        RECT  12.630 4.640 27.530 5.440 ;
        RECT  12.230 4.480 12.630 5.440 ;
        RECT  9.270 4.640 12.230 5.440 ;
        RECT  8.870 4.480 9.270 5.440 ;
        RECT  6.350 4.640 8.870 5.440 ;
        RECT  5.950 4.480 6.350 5.440 ;
        RECT  2.510 4.640 5.950 5.440 ;
        RECT  2.110 4.080 2.510 5.440 ;
        RECT  1.280 4.640 2.110 5.440 ;
        RECT  0.880 4.060 1.280 5.440 ;
        RECT  0.000 4.640 0.880 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  34.690 -0.400 35.640 0.400 ;
        RECT  34.290 -0.400 34.690 0.610 ;
        RECT  33.180 -0.400 34.290 0.400 ;
        RECT  32.940 -0.400 33.180 1.460 ;
        RECT  30.070 -0.400 32.940 0.400 ;
        RECT  29.670 -0.400 30.070 0.560 ;
        RECT  27.350 -0.400 29.670 0.400 ;
        RECT  26.950 -0.400 27.350 0.560 ;
        RECT  12.990 -0.400 26.950 0.400 ;
        RECT  12.590 -0.400 12.990 0.980 ;
        RECT  9.690 -0.400 12.590 0.400 ;
        RECT  9.290 -0.400 9.690 0.840 ;
        RECT  8.110 -0.400 9.290 0.400 ;
        RECT  7.710 -0.400 8.110 0.560 ;
        RECT  2.630 -0.400 7.710 0.400 ;
        RECT  2.230 -0.400 2.630 0.560 ;
        RECT  1.280 -0.400 2.230 0.400 ;
        RECT  0.880 -0.400 1.280 1.560 ;
        RECT  0.000 -0.400 0.880 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  34.740 2.030 34.960 2.430 ;
        RECT  34.500 2.030 34.740 3.600 ;
        RECT  33.340 3.360 34.500 3.600 ;
        RECT  33.820 1.340 34.060 3.120 ;
        RECT  33.660 1.340 33.820 1.580 ;
        RECT  32.860 2.880 33.820 3.120 ;
        RECT  33.100 3.360 33.340 4.370 ;
        RECT  31.260 4.130 33.100 4.370 ;
        RECT  32.700 2.040 32.870 2.280 ;
        RECT  32.620 2.880 32.860 3.890 ;
        RECT  32.460 0.800 32.700 2.280 ;
        RECT  31.740 3.650 32.620 3.890 ;
        RECT  24.490 0.800 32.460 1.040 ;
        RECT  32.220 3.170 32.380 3.410 ;
        RECT  31.980 1.370 32.220 3.410 ;
        RECT  31.500 2.140 31.740 3.890 ;
        RECT  31.260 1.350 31.580 1.750 ;
        RECT  31.020 1.350 31.260 4.370 ;
        RECT  30.540 1.330 30.780 4.220 ;
        RECT  30.060 1.280 30.300 2.700 ;
        RECT  25.770 1.280 30.060 1.520 ;
        RECT  29.180 1.760 29.420 4.270 ;
        RECT  28.880 1.760 29.180 2.000 ;
        RECT  29.020 3.370 29.180 4.270 ;
        RECT  27.290 3.600 29.020 3.840 ;
        RECT  27.040 3.100 28.570 3.340 ;
        RECT  27.040 1.760 28.140 2.000 ;
        RECT  27.050 3.600 27.290 4.400 ;
        RECT  23.610 4.160 27.050 4.400 ;
        RECT  26.810 1.760 27.040 3.340 ;
        RECT  26.800 1.760 26.810 3.920 ;
        RECT  26.570 2.350 26.800 3.920 ;
        RECT  24.970 3.680 26.570 3.920 ;
        RECT  26.330 1.760 26.560 2.000 ;
        RECT  26.090 1.760 26.330 3.440 ;
        RECT  25.930 3.200 26.090 3.440 ;
        RECT  25.690 1.280 25.770 1.840 ;
        RECT  25.450 1.280 25.690 3.440 ;
        RECT  25.370 1.280 25.450 1.840 ;
        RECT  25.210 3.200 25.450 3.440 ;
        RECT  24.730 1.440 24.970 3.920 ;
        RECT  24.450 3.440 24.730 3.840 ;
        RECT  24.250 0.800 24.490 1.970 ;
        RECT  19.660 1.730 24.250 1.970 ;
        RECT  23.770 0.740 24.010 1.140 ;
        RECT  19.450 0.740 23.770 0.980 ;
        RECT  23.370 2.930 23.610 4.400 ;
        RECT  20.880 2.930 23.370 3.170 ;
        RECT  19.150 1.250 23.330 1.490 ;
        RECT  19.420 1.730 19.660 3.920 ;
        RECT  18.540 3.680 19.420 3.920 ;
        RECT  19.020 3.200 19.180 3.440 ;
        RECT  18.910 0.640 19.150 1.490 ;
        RECT  18.780 2.160 19.020 3.440 ;
        RECT  13.470 0.640 18.910 0.880 ;
        RECT  18.670 2.160 18.780 2.400 ;
        RECT  18.430 1.120 18.670 2.400 ;
        RECT  18.300 2.670 18.540 3.920 ;
        RECT  13.950 1.120 18.430 1.360 ;
        RECT  18.190 2.670 18.300 2.910 ;
        RECT  17.950 1.600 18.190 2.910 ;
        RECT  15.070 1.600 17.950 1.840 ;
        RECT  17.020 3.750 17.420 4.400 ;
        RECT  16.140 4.160 17.020 4.400 ;
        RECT  16.770 2.080 16.970 2.320 ;
        RECT  16.530 2.080 16.770 2.880 ;
        RECT  16.140 2.640 16.530 2.880 ;
        RECT  15.550 2.080 16.250 2.320 ;
        RECT  15.900 2.640 16.140 4.400 ;
        RECT  13.110 4.160 15.900 4.400 ;
        RECT  15.550 3.040 15.660 3.920 ;
        RECT  15.420 2.080 15.550 3.920 ;
        RECT  15.310 2.080 15.420 3.280 ;
        RECT  13.590 3.680 15.420 3.920 ;
        RECT  14.990 1.600 15.070 2.820 ;
        RECT  14.830 1.600 14.990 3.440 ;
        RECT  14.750 2.580 14.830 3.440 ;
        RECT  14.550 3.200 14.750 3.440 ;
        RECT  14.510 1.600 14.590 1.840 ;
        RECT  14.270 1.600 14.510 2.940 ;
        RECT  14.190 1.600 14.270 1.840 ;
        RECT  14.230 2.700 14.270 2.940 ;
        RECT  13.990 2.700 14.230 3.440 ;
        RECT  12.930 2.180 14.030 2.420 ;
        RECT  13.830 3.200 13.990 3.440 ;
        RECT  13.710 1.120 13.950 1.940 ;
        RECT  11.850 1.700 13.710 1.940 ;
        RECT  13.350 3.520 13.590 3.920 ;
        RECT  13.230 0.640 13.470 1.460 ;
        RECT  12.930 3.520 13.350 3.760 ;
        RECT  10.760 1.220 13.230 1.460 ;
        RECT  12.870 4.000 13.110 4.400 ;
        RECT  12.690 2.180 12.930 3.760 ;
        RECT  11.990 4.000 12.870 4.240 ;
        RECT  12.530 2.640 12.690 3.760 ;
        RECT  11.510 3.520 12.530 3.760 ;
        RECT  10.170 0.740 12.350 0.980 ;
        RECT  11.750 4.000 11.990 4.400 ;
        RECT  11.610 1.700 11.850 3.280 ;
        RECT  9.780 4.160 11.750 4.400 ;
        RECT  11.450 3.040 11.610 3.280 ;
        RECT  11.270 3.520 11.510 3.920 ;
        RECT  10.380 3.680 11.270 3.920 ;
        RECT  10.520 1.220 10.760 1.820 ;
        RECT  10.380 2.060 10.550 2.300 ;
        RECT  6.980 1.580 10.520 1.820 ;
        RECT  10.140 2.060 10.380 3.920 ;
        RECT  9.930 0.740 10.170 1.340 ;
        RECT  9.660 3.340 10.140 3.740 ;
        RECT  7.460 1.100 9.930 1.340 ;
        RECT  9.540 4.000 9.780 4.400 ;
        RECT  3.220 4.000 9.540 4.240 ;
        RECT  8.840 2.060 9.080 3.740 ;
        RECT  8.180 2.060 8.840 2.460 ;
        RECT  4.060 3.500 8.840 3.740 ;
        RECT  8.080 2.720 8.480 3.260 ;
        RECT  6.490 3.020 8.080 3.260 ;
        RECT  7.220 0.640 7.460 1.340 ;
        RECT  6.970 2.540 7.300 2.780 ;
        RECT  6.280 0.640 7.220 0.880 ;
        RECT  6.970 1.160 6.980 1.820 ;
        RECT  6.730 1.160 6.970 2.780 ;
        RECT  6.580 1.160 6.730 1.400 ;
        RECT  6.280 1.710 6.490 3.260 ;
        RECT  6.250 0.640 6.280 3.260 ;
        RECT  6.040 0.640 6.250 1.950 ;
        RECT  5.140 3.020 5.560 3.260 ;
        RECT  5.140 1.380 5.470 1.780 ;
        RECT  4.900 1.380 5.140 3.260 ;
        RECT  4.550 0.660 4.950 1.060 ;
        RECT  4.780 2.030 4.900 2.430 ;
        RECT  4.540 2.750 4.590 3.150 ;
        RECT  4.540 0.820 4.550 1.060 ;
        RECT  4.300 0.820 4.540 3.150 ;
        RECT  2.000 0.820 4.300 1.060 ;
        RECT  3.820 1.380 4.060 3.740 ;
        RECT  3.550 2.840 3.820 3.740 ;
        RECT  3.260 1.380 3.420 1.780 ;
        RECT  3.020 1.380 3.260 3.120 ;
        RECT  2.980 3.570 3.220 4.240 ;
        RECT  2.830 2.720 3.020 3.120 ;
        RECT  0.480 3.570 2.980 3.810 ;
        RECT  2.350 2.070 2.750 2.470 ;
        RECT  2.000 2.110 2.350 2.460 ;
        RECT  1.760 0.820 2.000 3.120 ;
        RECT  1.600 1.420 1.760 1.820 ;
        RECT  1.600 2.720 1.760 3.120 ;
        RECT  0.480 0.900 0.560 1.800 ;
        RECT  0.240 0.900 0.480 4.160 ;
        RECT  0.160 0.900 0.240 1.800 ;
    END
END AFCSHCONX2

MACRO AFCSHCINX4
    CLASS CORE ;
    FOREIGN AFCSHCINX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 37.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  37.420 0.720 37.460 1.840 ;
        RECT  37.420 2.640 37.460 4.120 ;
        RECT  37.180 0.720 37.420 4.120 ;
        RECT  37.170 0.720 37.180 1.840 ;
        RECT  37.060 2.380 37.180 4.120 ;
        RECT  37.060 0.720 37.170 1.620 ;
        RECT  36.410 2.380 37.060 3.780 ;
        END
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  35.090 0.700 35.980 1.070 ;
        END
    END CS
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  22.650 2.220 25.320 2.460 ;
        RECT  22.650 3.660 25.320 3.900 ;
        RECT  22.330 2.220 22.650 2.660 ;
        RECT  22.330 3.500 22.650 3.900 ;
        RECT  21.890 2.220 22.330 3.900 ;
        RECT  21.790 2.220 21.890 2.460 ;
        RECT  21.790 3.660 21.890 3.900 ;
        END
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.010 2.220 21.090 2.460 ;
        RECT  21.010 3.660 21.090 3.900 ;
        RECT  20.570 2.220 21.010 3.900 ;
        RECT  20.250 2.220 20.570 2.660 ;
        RECT  20.250 3.500 20.570 3.900 ;
        RECT  17.560 2.220 20.250 2.460 ;
        RECT  17.560 3.660 20.250 3.900 ;
        END
    END CO0
    PIN CI1N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  30.560 2.270 31.200 2.720 ;
        END
    END CI1N
    PIN CI0N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  11.700 2.360 12.430 2.970 ;
        END
    END CI0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.690 2.760 9.700 3.760 ;
        RECT  9.360 2.380 9.690 3.760 ;
        RECT  8.000 3.520 9.360 3.760 ;
        RECT  8.270 1.910 8.510 2.360 ;
        RECT  8.000 2.120 8.270 2.360 ;
        RECT  7.760 2.120 8.000 3.760 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.370 1.810 1.870 2.660 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  36.670 4.640 37.620 5.440 ;
        RECT  36.270 4.020 36.670 5.440 ;
        RECT  35.730 4.640 36.270 5.440 ;
        RECT  35.330 3.770 35.730 5.440 ;
        RECT  31.810 4.640 35.330 5.440 ;
        RECT  31.410 3.370 31.810 5.440 ;
        RECT  30.090 4.640 31.410 5.440 ;
        RECT  28.690 4.370 30.090 5.440 ;
        RECT  14.160 4.640 28.690 5.440 ;
        RECT  12.760 4.480 14.160 5.440 ;
        RECT  11.260 4.640 12.760 5.440 ;
        RECT  10.860 4.480 11.260 5.440 ;
        RECT  9.960 4.640 10.860 5.440 ;
        RECT  9.560 4.480 9.960 5.440 ;
        RECT  2.260 4.640 9.560 5.440 ;
        RECT  1.310 4.360 2.260 5.440 ;
        RECT  0.000 4.640 1.310 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  36.670 -0.400 37.620 0.400 ;
        RECT  36.270 -0.400 36.670 1.370 ;
        RECT  34.850 -0.400 36.270 0.400 ;
        RECT  34.610 -0.400 34.850 1.780 ;
        RECT  31.740 -0.400 34.610 0.400 ;
        RECT  31.340 -0.400 31.740 0.560 ;
        RECT  30.130 -0.400 31.340 0.400 ;
        RECT  28.230 -0.400 30.130 0.560 ;
        RECT  11.330 -0.400 28.230 0.400 ;
        RECT  10.930 -0.400 11.330 0.900 ;
        RECT  10.000 -0.400 10.930 0.400 ;
        RECT  9.600 -0.400 10.000 0.900 ;
        RECT  2.360 -0.400 9.600 0.400 ;
        RECT  0.960 -0.400 2.360 0.560 ;
        RECT  0.000 -0.400 0.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  36.170 1.890 36.930 2.130 ;
        RECT  35.930 1.890 36.170 3.530 ;
        RECT  35.090 3.290 35.930 3.530 ;
        RECT  35.360 2.810 35.690 3.050 ;
        RECT  35.360 1.380 35.680 1.620 ;
        RECT  35.120 1.380 35.360 3.050 ;
        RECT  34.610 2.810 35.120 3.050 ;
        RECT  34.850 3.290 35.090 4.400 ;
        RECT  33.170 4.160 34.850 4.400 ;
        RECT  34.370 2.810 34.610 3.920 ;
        RECT  34.370 2.020 34.580 2.260 ;
        RECT  34.130 0.800 34.370 2.260 ;
        RECT  33.650 3.680 34.370 3.920 ;
        RECT  25.710 0.800 34.130 1.040 ;
        RECT  33.890 2.500 34.130 3.440 ;
        RECT  33.650 1.350 33.890 2.740 ;
        RECT  33.410 2.980 33.650 3.920 ;
        RECT  33.170 2.140 33.410 3.220 ;
        RECT  32.930 1.350 33.250 1.750 ;
        RECT  32.930 3.500 33.170 4.400 ;
        RECT  32.690 1.350 32.930 4.400 ;
        RECT  32.210 1.350 32.450 4.010 ;
        RECT  31.900 2.360 31.960 2.760 ;
        RECT  31.660 1.280 31.900 2.760 ;
        RECT  27.120 1.280 31.660 1.520 ;
        RECT  30.690 2.980 31.090 4.380 ;
        RECT  30.210 1.760 30.950 2.000 ;
        RECT  30.210 3.570 30.690 3.910 ;
        RECT  29.970 1.760 30.210 3.910 ;
        RECT  26.400 3.670 29.970 3.910 ;
        RECT  29.420 2.980 29.720 3.380 ;
        RECT  29.420 1.760 29.580 2.000 ;
        RECT  29.180 1.760 29.420 3.380 ;
        RECT  28.260 2.350 29.180 2.750 ;
        RECT  28.020 2.990 28.260 3.390 ;
        RECT  15.170 4.160 28.030 4.400 ;
        RECT  27.780 1.760 28.020 3.390 ;
        RECT  27.440 1.760 27.780 2.000 ;
        RECT  27.140 2.990 27.540 3.390 ;
        RECT  27.120 2.990 27.140 3.230 ;
        RECT  26.880 1.280 27.120 3.230 ;
        RECT  26.720 1.550 26.880 1.950 ;
        RECT  26.160 1.610 26.400 3.910 ;
        RECT  26.000 1.610 26.160 3.180 ;
        RECT  22.690 2.940 26.000 3.180 ;
        RECT  25.470 0.800 25.710 1.980 ;
        RECT  17.520 1.740 25.470 1.980 ;
        RECT  21.820 1.250 25.190 1.490 ;
        RECT  21.580 0.640 21.820 1.490 ;
        RECT  11.810 0.640 21.580 0.880 ;
        RECT  18.130 1.250 21.100 1.490 ;
        RECT  17.040 2.940 20.160 3.180 ;
        RECT  17.810 1.120 18.130 1.490 ;
        RECT  12.290 1.120 17.810 1.360 ;
        RECT  17.280 1.600 17.520 1.980 ;
        RECT  16.250 1.600 17.280 1.840 ;
        RECT  16.800 2.080 17.040 3.760 ;
        RECT  16.640 2.080 16.800 2.320 ;
        RECT  16.530 3.520 16.800 3.760 ;
        RECT  16.130 3.520 16.530 3.910 ;
        RECT  16.170 1.600 16.250 2.000 ;
        RECT  15.930 1.600 16.170 3.280 ;
        RECT  12.910 3.520 16.130 3.760 ;
        RECT  15.850 1.600 15.930 2.000 ;
        RECT  15.340 3.040 15.930 3.280 ;
        RECT  15.130 1.660 15.530 2.060 ;
        RECT  14.850 4.000 15.170 4.400 ;
        RECT  15.100 1.820 15.130 2.060 ;
        RECT  14.860 1.820 15.100 3.280 ;
        RECT  14.620 3.040 14.860 3.280 ;
        RECT  7.510 4.000 14.850 4.240 ;
        RECT  14.220 2.350 14.620 2.750 ;
        RECT  13.980 1.640 14.220 3.270 ;
        RECT  13.820 1.640 13.980 2.040 ;
        RECT  13.240 3.030 13.980 3.270 ;
        RECT  12.670 1.640 12.910 3.760 ;
        RECT  12.530 1.640 12.670 2.040 ;
        RECT  11.650 3.360 12.670 3.760 ;
        RECT  12.050 1.120 12.290 1.860 ;
        RECT  10.910 1.620 12.050 1.860 ;
        RECT  11.570 0.640 11.810 1.380 ;
        RECT  9.130 1.140 11.570 1.380 ;
        RECT  10.670 1.620 10.910 3.640 ;
        RECT  10.420 1.620 10.670 2.020 ;
        RECT  10.350 3.240 10.670 3.640 ;
        RECT  10.180 2.260 10.400 2.660 ;
        RECT  9.940 1.620 10.180 2.660 ;
        RECT  9.100 1.620 9.940 1.860 ;
        RECT  8.890 0.640 9.130 1.380 ;
        RECT  8.860 1.620 9.100 3.240 ;
        RECT  7.500 0.640 8.890 0.880 ;
        RECT  8.480 3.000 8.860 3.240 ;
        RECT  7.980 1.230 8.620 1.630 ;
        RECT  8.240 2.670 8.480 3.240 ;
        RECT  7.740 1.230 7.980 1.840 ;
        RECT  6.780 1.600 7.740 1.840 ;
        RECT  7.270 2.940 7.510 4.240 ;
        RECT  7.260 0.640 7.500 1.360 ;
        RECT  7.020 2.140 7.420 2.700 ;
        RECT  6.410 2.940 7.270 3.180 ;
        RECT  6.300 1.120 7.260 1.360 ;
        RECT  5.590 0.640 7.020 0.880 ;
        RECT  5.590 2.460 7.020 2.700 ;
        RECT  6.930 3.580 7.020 3.980 ;
        RECT  6.690 3.580 6.930 4.360 ;
        RECT  6.540 1.600 6.780 2.200 ;
        RECT  3.890 4.120 6.690 4.360 ;
        RECT  4.190 1.960 6.540 2.200 ;
        RECT  6.170 2.940 6.410 3.560 ;
        RECT  6.060 1.120 6.300 1.720 ;
        RECT  5.590 3.320 6.170 3.560 ;
        RECT  3.250 1.480 6.060 1.720 ;
        RECT  5.350 0.640 5.590 1.240 ;
        RECT  5.350 2.460 5.590 3.000 ;
        RECT  4.190 3.320 5.590 3.720 ;
        RECT  4.190 0.800 5.350 1.240 ;
        RECT  4.190 2.600 5.350 3.000 ;
        RECT  0.560 0.800 4.190 1.040 ;
        RECT  3.920 2.760 4.190 3.000 ;
        RECT  3.680 2.760 3.920 3.620 ;
        RECT  3.650 3.870 3.890 4.360 ;
        RECT  1.860 3.380 3.680 3.620 ;
        RECT  0.560 3.870 3.650 4.110 ;
        RECT  3.010 1.320 3.250 3.140 ;
        RECT  2.760 1.320 3.010 1.720 ;
        RECT  2.760 2.740 3.010 3.140 ;
        RECT  2.510 2.040 2.770 2.440 ;
        RECT  2.270 1.280 2.510 2.440 ;
        RECT  1.040 1.280 2.270 1.520 ;
        RECT  1.460 3.050 1.860 3.620 ;
        RECT  1.040 3.050 1.460 3.290 ;
        RECT  0.800 1.280 1.040 3.290 ;
        RECT  0.630 2.080 0.800 2.480 ;
        RECT  0.370 0.720 0.560 1.620 ;
        RECT  0.370 2.820 0.560 4.220 ;
        RECT  0.130 0.720 0.370 4.220 ;
    END
END AFCSHCINX4

MACRO AFCSHCINX2
    CLASS CORE ;
    FOREIGN AFCSHCINX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AFCSHCINX4 ;
    SIZE 36.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  36.760 0.720 36.800 1.840 ;
        RECT  36.760 2.640 36.800 4.120 ;
        RECT  36.520 0.720 36.760 4.120 ;
        RECT  36.510 0.720 36.520 1.840 ;
        RECT  36.400 2.380 36.520 4.120 ;
        RECT  36.400 0.720 36.510 1.620 ;
        RECT  35.750 2.380 36.400 3.780 ;
        END
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  34.430 0.700 35.320 1.070 ;
        END
    END CS
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  22.650 3.660 25.450 3.900 ;
        RECT  22.330 2.140 25.280 2.380 ;
        RECT  22.330 3.500 22.650 3.900 ;
        RECT  21.890 2.140 22.330 3.900 ;
        RECT  21.790 2.140 21.890 2.380 ;
        END
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.010 2.140 21.090 2.380 ;
        RECT  20.570 2.140 21.010 3.890 ;
        RECT  17.560 2.140 20.570 2.380 ;
        RECT  20.240 3.500 20.570 3.890 ;
        RECT  17.590 3.650 20.240 3.890 ;
        END
    END CO0
    PIN CI1N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  29.640 2.270 30.250 2.720 ;
        END
    END CI1N
    PIN CI0N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  11.700 2.360 12.430 2.970 ;
        END
    END CI0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.690 2.760 9.700 3.760 ;
        RECT  9.360 2.380 9.690 3.760 ;
        RECT  8.000 3.520 9.360 3.760 ;
        RECT  8.270 1.910 8.510 2.360 ;
        RECT  8.000 2.120 8.270 2.360 ;
        RECT  7.760 2.120 8.000 3.760 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.370 1.810 1.870 2.660 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  36.010 4.640 36.960 5.440 ;
        RECT  35.610 4.020 36.010 5.440 ;
        RECT  35.070 4.640 35.610 5.440 ;
        RECT  34.670 3.770 35.070 5.440 ;
        RECT  31.150 4.640 34.670 5.440 ;
        RECT  30.750 3.500 31.150 5.440 ;
        RECT  29.590 4.640 30.750 5.440 ;
        RECT  28.690 4.370 29.590 5.440 ;
        RECT  13.970 4.640 28.690 5.440 ;
        RECT  12.570 4.480 13.970 5.440 ;
        RECT  11.490 4.640 12.570 5.440 ;
        RECT  11.090 4.480 11.490 5.440 ;
        RECT  9.960 4.640 11.090 5.440 ;
        RECT  9.560 4.480 9.960 5.440 ;
        RECT  2.260 4.640 9.560 5.440 ;
        RECT  1.310 4.360 2.260 5.440 ;
        RECT  0.000 4.640 1.310 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  36.010 -0.400 36.960 0.400 ;
        RECT  35.610 -0.400 36.010 1.370 ;
        RECT  34.190 -0.400 35.610 0.400 ;
        RECT  33.950 -0.400 34.190 1.780 ;
        RECT  31.080 -0.400 33.950 0.400 ;
        RECT  30.680 -0.400 31.080 0.560 ;
        RECT  29.100 -0.400 30.680 0.400 ;
        RECT  28.200 -0.400 29.100 0.560 ;
        RECT  11.330 -0.400 28.200 0.400 ;
        RECT  10.930 -0.400 11.330 0.900 ;
        RECT  10.000 -0.400 10.930 0.400 ;
        RECT  9.600 -0.400 10.000 0.900 ;
        RECT  2.360 -0.400 9.600 0.400 ;
        RECT  0.960 -0.400 2.360 0.560 ;
        RECT  0.000 -0.400 0.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  35.510 1.890 36.270 2.130 ;
        RECT  35.270 1.890 35.510 3.530 ;
        RECT  34.430 3.290 35.270 3.530 ;
        RECT  34.700 2.810 35.030 3.050 ;
        RECT  34.700 1.380 35.020 1.620 ;
        RECT  34.460 1.380 34.700 3.050 ;
        RECT  33.950 2.810 34.460 3.050 ;
        RECT  34.190 3.290 34.430 4.400 ;
        RECT  32.510 4.160 34.190 4.400 ;
        RECT  33.710 2.810 33.950 3.920 ;
        RECT  33.710 2.020 33.920 2.260 ;
        RECT  33.470 0.800 33.710 2.260 ;
        RECT  32.990 3.680 33.710 3.920 ;
        RECT  25.760 0.800 33.470 1.040 ;
        RECT  33.230 2.500 33.470 3.440 ;
        RECT  32.990 1.350 33.230 2.740 ;
        RECT  32.750 2.980 32.990 3.920 ;
        RECT  32.510 2.140 32.750 3.220 ;
        RECT  32.270 1.350 32.590 1.750 ;
        RECT  32.270 3.460 32.510 4.400 ;
        RECT  32.030 1.350 32.270 4.400 ;
        RECT  31.550 1.350 31.790 4.170 ;
        RECT  31.240 2.360 31.300 2.760 ;
        RECT  31.000 1.280 31.240 2.760 ;
        RECT  27.120 1.280 31.000 1.520 ;
        RECT  30.520 1.760 30.760 3.220 ;
        RECT  29.890 1.760 30.520 2.000 ;
        RECT  30.430 2.980 30.520 3.220 ;
        RECT  30.030 2.980 30.430 4.380 ;
        RECT  26.400 3.670 30.030 3.910 ;
        RECT  29.320 3.060 29.630 3.300 ;
        RECT  29.320 1.760 29.480 2.000 ;
        RECT  29.080 1.760 29.320 3.300 ;
        RECT  28.180 2.350 29.080 2.750 ;
        RECT  27.940 2.990 28.260 3.390 ;
        RECT  15.170 4.160 28.030 4.400 ;
        RECT  27.700 1.760 27.940 3.390 ;
        RECT  27.440 1.760 27.700 2.000 ;
        RECT  27.220 2.990 27.460 3.390 ;
        RECT  27.120 2.990 27.220 3.230 ;
        RECT  26.880 1.280 27.120 3.230 ;
        RECT  26.720 1.550 26.880 1.950 ;
        RECT  26.160 1.530 26.400 3.910 ;
        RECT  26.000 1.530 26.160 3.170 ;
        RECT  25.450 2.930 26.000 3.170 ;
        RECT  25.520 0.800 25.760 1.840 ;
        RECT  16.170 1.600 25.520 1.840 ;
        RECT  24.890 2.930 25.450 3.180 ;
        RECT  21.820 1.120 25.280 1.360 ;
        RECT  22.690 2.930 24.890 3.170 ;
        RECT  21.580 0.640 21.820 1.360 ;
        RECT  11.810 0.640 21.580 0.880 ;
        RECT  12.290 1.120 21.100 1.360 ;
        RECT  16.650 2.930 20.140 3.170 ;
        RECT  16.650 2.080 17.040 2.320 ;
        RECT  16.530 2.080 16.650 3.820 ;
        RECT  16.410 2.080 16.530 3.910 ;
        RECT  16.130 3.520 16.410 3.910 ;
        RECT  15.930 1.600 16.170 3.280 ;
        RECT  12.910 3.520 16.130 3.760 ;
        RECT  15.340 3.040 15.930 3.280 ;
        RECT  15.130 1.660 15.530 2.060 ;
        RECT  14.850 4.000 15.170 4.400 ;
        RECT  15.100 1.820 15.130 2.060 ;
        RECT  14.860 1.820 15.100 3.280 ;
        RECT  14.620 3.040 14.860 3.280 ;
        RECT  7.510 4.000 14.850 4.240 ;
        RECT  13.710 2.350 14.620 2.750 ;
        RECT  13.470 1.640 13.710 3.270 ;
        RECT  13.310 1.640 13.470 2.040 ;
        RECT  13.240 3.030 13.470 3.270 ;
        RECT  12.670 1.640 12.910 3.760 ;
        RECT  12.530 1.640 12.670 2.040 ;
        RECT  11.690 3.360 12.670 3.760 ;
        RECT  12.050 1.120 12.290 1.860 ;
        RECT  10.910 1.620 12.050 1.860 ;
        RECT  11.570 0.640 11.810 1.380 ;
        RECT  9.130 1.140 11.570 1.380 ;
        RECT  10.670 1.620 10.910 3.640 ;
        RECT  10.420 1.620 10.670 2.020 ;
        RECT  10.350 3.240 10.670 3.640 ;
        RECT  10.180 2.260 10.400 2.660 ;
        RECT  9.940 1.620 10.180 2.660 ;
        RECT  9.100 1.620 9.940 1.860 ;
        RECT  8.890 0.640 9.130 1.380 ;
        RECT  8.860 1.620 9.100 3.240 ;
        RECT  7.500 0.640 8.890 0.880 ;
        RECT  8.480 3.000 8.860 3.240 ;
        RECT  7.980 1.230 8.620 1.630 ;
        RECT  8.240 2.670 8.480 3.240 ;
        RECT  7.740 1.230 7.980 1.840 ;
        RECT  6.550 1.600 7.740 1.840 ;
        RECT  7.270 2.940 7.510 4.240 ;
        RECT  7.260 0.640 7.500 1.360 ;
        RECT  7.020 2.140 7.420 2.700 ;
        RECT  6.410 2.940 7.270 3.180 ;
        RECT  6.070 1.120 7.260 1.360 ;
        RECT  5.590 0.640 7.020 0.880 ;
        RECT  5.640 2.460 7.020 2.700 ;
        RECT  6.930 3.580 7.020 3.980 ;
        RECT  6.690 3.580 6.930 4.360 ;
        RECT  3.890 4.120 6.690 4.360 ;
        RECT  6.310 1.600 6.550 2.200 ;
        RECT  6.170 2.940 6.410 3.560 ;
        RECT  4.190 1.960 6.310 2.200 ;
        RECT  5.610 3.320 6.170 3.560 ;
        RECT  5.830 1.120 6.070 1.720 ;
        RECT  3.250 1.480 5.830 1.720 ;
        RECT  5.400 2.460 5.640 3.000 ;
        RECT  4.210 3.320 5.610 3.720 ;
        RECT  5.350 0.640 5.590 1.240 ;
        RECT  4.240 2.600 5.400 3.000 ;
        RECT  4.190 0.800 5.350 1.240 ;
        RECT  3.920 2.760 4.240 3.000 ;
        RECT  0.560 0.800 4.190 1.040 ;
        RECT  3.680 2.760 3.920 3.620 ;
        RECT  3.650 3.870 3.890 4.360 ;
        RECT  1.860 3.380 3.680 3.620 ;
        RECT  0.560 3.870 3.650 4.110 ;
        RECT  3.010 1.320 3.250 3.140 ;
        RECT  2.760 1.320 3.010 1.720 ;
        RECT  2.760 2.740 3.010 3.140 ;
        RECT  2.510 2.040 2.770 2.440 ;
        RECT  2.270 1.280 2.510 2.440 ;
        RECT  1.130 1.280 2.270 1.520 ;
        RECT  1.460 3.050 1.860 3.620 ;
        RECT  1.130 3.050 1.460 3.290 ;
        RECT  0.890 1.280 1.130 3.290 ;
        RECT  0.630 2.080 0.890 2.480 ;
        RECT  0.370 0.720 0.560 1.620 ;
        RECT  0.370 2.820 0.560 4.220 ;
        RECT  0.130 0.720 0.370 4.220 ;
    END
END AFCSHCINX2

MACRO AHHCONX4
    CLASS CORE ;
    FOREIGN AHHCONX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.240 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.940 2.950 3.090 3.190 ;
        RECT  3.090 2.950 3.260 3.220 ;
        RECT  3.260 2.950 3.500 3.680 ;
        RECT  3.340 0.670 4.230 0.910 ;
        RECT  4.230 0.670 4.470 1.060 ;
        RECT  4.470 0.820 4.730 1.060 ;
        RECT  3.500 3.440 4.740 3.680 ;
        RECT  4.730 0.820 4.740 2.660 ;
        RECT  4.740 0.820 4.970 3.680 ;
        RECT  4.970 1.260 4.980 3.680 ;
        RECT  4.980 1.260 5.170 2.660 ;
        END
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  5.240 3.150 5.730 3.390 ;
        RECT  5.730 2.940 6.050 3.390 ;
        RECT  6.050 1.820 6.180 3.390 ;
        RECT  6.180 1.150 6.420 3.390 ;
        RECT  6.420 1.820 6.490 3.390 ;
        RECT  6.490 2.380 6.810 3.390 ;
        RECT  6.810 2.500 7.230 3.390 ;
        RECT  7.230 2.500 7.620 2.740 ;
        RECT  7.620 1.310 7.860 2.740 ;
        RECT  7.860 1.310 8.370 1.550 ;
        RECT  8.370 1.150 8.860 1.550 ;
        END
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.850 2.330 1.930 2.570 ;
        RECT  1.930 2.280 2.250 2.570 ;
        RECT  2.250 2.280 2.490 3.760 ;
        RECT  2.490 3.510 2.780 3.760 ;
        RECT  2.780 3.510 3.020 4.220 ;
        RECT  3.020 3.980 3.410 4.220 ;
        RECT  2.490 2.280 3.650 2.520 ;
        RECT  3.410 3.980 3.850 4.340 ;
        RECT  3.650 1.840 3.890 2.520 ;
        RECT  3.850 3.980 7.500 4.220 ;
        RECT  7.500 2.990 7.740 4.220 ;
        RECT  7.740 2.990 8.310 3.230 ;
        RECT  8.310 2.260 8.550 3.230 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.540 0.670 5.780 2.660 ;
        RECT  5.780 0.670 6.710 0.910 ;
        RECT  6.710 0.670 6.950 1.550 ;
        RECT  6.950 1.270 7.060 1.550 ;
        RECT  7.060 1.310 7.130 1.550 ;
        RECT  7.130 1.310 7.370 2.090 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.000 5.440 ;
        RECT  1.000 4.480 1.400 5.440 ;
        RECT  1.400 4.640 4.450 5.440 ;
        RECT  4.450 4.480 4.850 5.440 ;
        RECT  4.850 4.640 6.030 5.440 ;
        RECT  6.030 4.480 6.430 5.440 ;
        RECT  6.430 4.640 7.700 5.440 ;
        RECT  7.700 4.480 8.090 5.440 ;
        RECT  8.090 3.750 8.490 5.440 ;
        RECT  8.490 4.640 9.240 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.000 0.400 ;
        RECT  1.000 -0.400 1.400 0.560 ;
        RECT  1.400 -0.400 4.850 0.400 ;
        RECT  4.850 -0.400 5.250 0.560 ;
        RECT  5.250 -0.400 7.280 0.400 ;
        RECT  7.280 -0.400 7.680 0.850 ;
        RECT  7.680 -0.400 9.240 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.450 1.360 4.460 1.600 ;
        RECT  4.210 1.360 4.450 3.030 ;
        RECT  3.170 1.360 4.210 1.600 ;
        RECT  3.980 2.790 4.210 3.030 ;
        RECT  3.740 2.790 3.980 3.200 ;
        RECT  2.930 1.360 3.170 2.030 ;
        RECT  1.490 1.790 2.930 2.030 ;
        RECT  2.450 0.640 2.690 1.040 ;
        RECT  2.650 1.280 2.670 1.520 ;
        RECT  2.270 1.280 2.650 1.530 ;
        RECT  2.300 4.000 2.540 4.400 ;
        RECT  0.530 0.800 2.450 1.040 ;
        RECT  0.530 4.000 2.300 4.240 ;
        RECT  1.010 1.290 2.270 1.530 ;
        RECT  1.600 3.150 2.000 3.550 ;
        RECT  1.010 3.150 1.600 3.390 ;
        RECT  1.250 1.790 1.490 2.580 ;
        RECT  0.770 1.290 1.010 3.390 ;
        RECT  0.290 0.800 0.530 4.240 ;
    END
END AHHCONX4

MACRO AHHCONX2
    CLASS CORE ;
    FOREIGN AHHCONX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AHHCONX4 ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.950 3.100 3.210 ;
        RECT  3.100 2.840 3.340 3.200 ;
        RECT  3.420 1.170 3.660 1.580 ;
        RECT  3.340 2.840 4.110 3.080 ;
        RECT  3.660 1.340 4.110 1.580 ;
        RECT  4.110 1.340 4.350 3.080 ;
        END
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  5.240 3.080 6.070 3.320 ;
        RECT  6.070 1.280 6.100 3.320 ;
        RECT  6.100 1.120 6.310 3.320 ;
        RECT  6.310 1.120 6.500 1.540 ;
        RECT  6.500 1.260 7.150 1.540 ;
        END
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.850 2.330 2.250 2.570 ;
        RECT  2.250 2.330 2.490 3.760 ;
        RECT  2.490 3.510 2.870 3.760 ;
        RECT  2.870 3.510 3.110 4.040 ;
        RECT  3.110 3.700 3.190 4.040 ;
        RECT  3.190 3.800 3.410 4.040 ;
        RECT  2.490 2.330 3.410 2.570 ;
        RECT  3.410 2.080 3.630 2.570 ;
        RECT  3.410 3.800 3.850 4.340 ;
        RECT  3.630 1.840 3.870 2.570 ;
        RECT  3.850 3.800 6.550 4.040 ;
        RECT  6.550 2.250 6.790 4.040 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.070 1.820 5.830 2.310 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.000 5.440 ;
        RECT  1.000 4.480 1.400 5.440 ;
        RECT  1.400 4.640 4.450 5.440 ;
        RECT  4.450 4.480 4.850 5.440 ;
        RECT  4.850 4.640 6.030 5.440 ;
        RECT  6.030 4.480 6.430 5.440 ;
        RECT  6.430 4.640 7.920 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.000 0.400 ;
        RECT  1.000 -0.400 1.400 0.560 ;
        RECT  1.400 -0.400 4.850 0.400 ;
        RECT  4.850 -0.400 5.250 0.560 ;
        RECT  5.250 -0.400 7.350 0.400 ;
        RECT  7.350 -0.400 7.750 0.560 ;
        RECT  7.750 -0.400 7.920 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.610 0.800 4.830 3.560 ;
        RECT  4.590 0.690 4.610 3.560 ;
        RECT  4.370 0.690 4.590 1.040 ;
        RECT  3.660 3.320 4.590 3.560 ;
        RECT  3.170 0.690 4.370 0.930 ;
        RECT  2.930 0.690 3.170 2.030 ;
        RECT  1.490 1.790 2.930 2.030 ;
        RECT  2.450 0.640 2.690 1.040 ;
        RECT  2.650 1.280 2.670 1.520 ;
        RECT  2.270 1.280 2.650 1.530 ;
        RECT  0.530 4.000 2.620 4.240 ;
        RECT  0.530 0.800 2.450 1.040 ;
        RECT  1.010 1.290 2.270 1.530 ;
        RECT  1.600 3.150 2.000 3.550 ;
        RECT  1.010 3.150 1.600 3.390 ;
        RECT  1.250 1.790 1.490 2.580 ;
        RECT  0.770 1.290 1.010 3.390 ;
        RECT  0.290 0.800 0.530 4.240 ;
    END
END AHHCONX2

MACRO AHHCINX4
    CLASS CORE ;
    FOREIGN AHHCINX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.590 1.220 3.610 2.080 ;
        RECT  3.370 1.220 3.590 3.900 ;
        RECT  3.210 1.820 3.370 3.900 ;
        RECT  2.750 1.820 3.210 3.220 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.500 1.620 9.740 2.980 ;
        RECT  8.490 1.620 9.500 1.860 ;
        RECT  9.050 2.740 9.500 2.980 ;
        RECT  8.580 2.740 9.050 3.620 ;
        RECT  8.030 2.740 8.580 4.340 ;
        RECT  8.250 1.300 8.490 1.860 ;
        RECT  7.350 1.300 8.250 1.540 ;
        RECT  6.810 2.760 8.030 3.000 ;
        RECT  6.950 0.670 7.350 1.540 ;
        RECT  5.850 1.210 6.950 1.450 ;
        RECT  6.550 2.760 6.810 3.220 ;
        RECT  6.150 2.760 6.550 4.180 ;
        RECT  5.450 0.670 5.850 1.450 ;
        END
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.760 2.260 7.500 2.500 ;
        RECT  5.560 2.260 5.760 3.240 ;
        RECT  5.320 2.180 5.560 3.720 ;
        RECT  4.250 3.480 5.320 3.720 ;
        RECT  4.010 3.480 4.250 4.400 ;
        RECT  1.710 4.160 4.010 4.400 ;
        END
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.840 2.100 9.240 2.500 ;
        RECT  8.000 2.100 8.840 2.340 ;
        RECT  7.760 1.780 8.000 2.340 ;
        RECT  6.450 1.780 7.760 2.020 ;
        RECT  6.210 1.700 6.450 2.020 ;
        RECT  5.170 1.700 6.210 1.940 ;
        RECT  4.970 1.260 5.170 1.940 ;
        RECT  4.730 1.260 4.970 2.340 ;
        RECT  4.330 1.940 4.730 2.340 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  9.590 4.640 10.560 5.440 ;
        RECT  9.190 3.940 9.590 5.440 ;
        RECT  7.780 4.640 9.190 5.440 ;
        RECT  7.420 3.260 7.780 5.440 ;
        RECT  6.200 4.600 7.420 5.440 ;
        RECT  5.140 4.640 6.200 5.440 ;
        RECT  4.740 3.980 5.140 5.440 ;
        RECT  1.420 4.640 4.740 5.440 ;
        RECT  1.020 4.420 1.420 5.440 ;
        RECT  0.000 4.640 1.020 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  9.460 -0.400 10.560 0.400 ;
        RECT  8.570 -0.400 9.460 0.620 ;
        RECT  8.010 -0.400 8.570 1.060 ;
        RECT  6.570 -0.400 8.010 0.400 ;
        RECT  7.670 0.820 8.010 1.060 ;
        RECT  6.170 -0.400 6.570 0.940 ;
        RECT  5.130 -0.400 6.170 0.400 ;
        RECT  4.730 -0.400 5.130 0.940 ;
        RECT  1.940 -0.400 4.730 0.400 ;
        RECT  0.930 -0.400 1.940 0.560 ;
        RECT  0.000 -0.400 0.930 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.300 0.640 10.400 1.540 ;
        RECT  10.300 2.720 10.400 4.280 ;
        RECT  10.000 0.640 10.300 4.280 ;
        RECT  9.240 0.980 10.000 1.280 ;
        RECT  8.840 0.980 9.240 1.380 ;
        RECT  4.090 0.690 4.410 1.590 ;
        RECT  4.090 2.820 4.350 3.220 ;
        RECT  3.850 0.690 4.090 3.220 ;
        RECT  3.130 0.690 3.850 0.930 ;
        RECT  2.890 0.690 3.130 1.530 ;
        RECT  2.510 3.490 2.910 3.920 ;
        RECT  2.510 1.290 2.890 1.530 ;
        RECT  2.410 0.640 2.650 1.040 ;
        RECT  2.270 1.290 2.510 2.020 ;
        RECT  0.630 3.680 2.510 3.920 ;
        RECT  2.260 2.300 2.500 3.060 ;
        RECT  0.630 0.800 2.410 1.040 ;
        RECT  1.950 1.780 2.270 2.020 ;
        RECT  1.990 2.820 2.260 3.060 ;
        RECT  1.440 1.280 2.010 1.520 ;
        RECT  1.570 2.820 1.990 3.440 ;
        RECT  1.710 1.780 1.950 2.400 ;
        RECT  1.400 2.160 1.710 2.400 ;
        RECT  0.920 2.820 1.570 3.060 ;
        RECT  1.200 1.280 1.440 1.910 ;
        RECT  1.160 2.160 1.400 2.560 ;
        RECT  0.920 1.670 1.200 1.910 ;
        RECT  0.680 1.670 0.920 3.060 ;
        RECT  0.440 0.660 0.630 1.430 ;
        RECT  0.440 3.340 0.630 4.240 ;
        RECT  0.200 0.660 0.440 4.240 ;
    END
END AHHCINX4

MACRO AHHCINX2
    CLASS CORE ;
    FOREIGN AHHCINX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AHHCINX4 ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.370 1.220 3.610 3.770 ;
        RECT  3.250 2.860 3.370 3.770 ;
        RECT  2.750 2.940 3.250 3.220 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.230 1.350 6.470 3.220 ;
        RECT  5.850 1.350 6.230 1.590 ;
        RECT  5.450 0.640 5.850 1.590 ;
        END
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.190 2.280 7.430 4.240 ;
        RECT  5.510 4.000 7.190 4.240 ;
        RECT  5.110 2.340 5.510 4.240 ;
        RECT  4.410 4.000 5.110 4.240 ;
        RECT  4.170 4.000 4.410 4.400 ;
        RECT  3.410 4.060 4.170 4.400 ;
        RECT  1.650 4.160 3.410 4.400 ;
        END
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.500 1.600 7.900 2.040 ;
        RECT  6.950 1.800 7.500 2.040 ;
        RECT  6.710 1.800 6.950 3.740 ;
        RECT  5.990 3.500 6.710 3.740 ;
        RECT  5.750 1.830 5.990 3.740 ;
        RECT  5.080 1.830 5.750 2.070 ;
        RECT  4.830 1.830 5.080 2.090 ;
        RECT  4.430 1.830 4.830 2.580 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  7.810 4.640 8.580 5.440 ;
        RECT  7.410 4.480 7.810 5.440 ;
        RECT  6.760 4.640 7.410 5.440 ;
        RECT  5.820 4.600 6.760 5.440 ;
        RECT  5.140 4.640 5.820 5.440 ;
        RECT  4.740 4.480 5.140 5.440 ;
        RECT  1.420 4.640 4.740 5.440 ;
        RECT  1.020 4.480 1.420 5.440 ;
        RECT  0.000 4.640 1.020 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  7.180 -0.400 8.580 0.400 ;
        RECT  6.570 -0.400 7.180 0.600 ;
        RECT  6.170 -0.400 6.570 1.080 ;
        RECT  5.130 -0.400 6.170 0.400 ;
        RECT  4.730 -0.400 5.130 1.440 ;
        RECT  1.940 -0.400 4.730 0.400 ;
        RECT  0.930 -0.400 1.940 0.560 ;
        RECT  0.000 -0.400 0.930 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  8.380 3.020 8.420 3.420 ;
        RECT  8.250 1.120 8.380 3.420 ;
        RECT  8.140 0.840 8.250 3.420 ;
        RECT  7.850 0.840 8.140 1.360 ;
        RECT  8.020 3.020 8.140 3.420 ;
        RECT  7.180 1.120 7.850 1.360 ;
        RECT  6.810 1.120 7.180 1.560 ;
        RECT  6.780 1.320 6.810 1.560 ;
        RECT  4.110 0.660 4.410 1.560 ;
        RECT  4.110 2.860 4.350 3.760 ;
        RECT  4.010 0.660 4.110 3.760 ;
        RECT  3.870 0.710 4.010 3.760 ;
        RECT  3.130 0.710 3.870 0.950 ;
        RECT  2.890 0.710 3.130 2.090 ;
        RECT  2.510 3.470 2.910 3.920 ;
        RECT  1.940 1.850 2.890 2.090 ;
        RECT  2.410 0.650 2.650 1.550 ;
        RECT  2.420 2.380 2.580 2.620 ;
        RECT  0.630 3.680 2.510 3.920 ;
        RECT  2.180 2.380 2.420 3.060 ;
        RECT  0.630 0.800 2.410 1.040 ;
        RECT  1.990 2.820 2.180 3.060 ;
        RECT  1.440 1.280 2.010 1.520 ;
        RECT  1.590 2.820 1.990 3.440 ;
        RECT  1.700 1.850 1.940 2.400 ;
        RECT  1.400 2.160 1.700 2.400 ;
        RECT  0.920 2.820 1.590 3.060 ;
        RECT  1.200 1.280 1.440 1.910 ;
        RECT  1.160 2.160 1.400 2.560 ;
        RECT  0.920 1.670 1.200 1.910 ;
        RECT  0.680 1.670 0.920 3.060 ;
        RECT  0.440 0.660 0.630 1.430 ;
        RECT  0.440 3.390 0.630 4.290 ;
        RECT  0.200 0.660 0.440 4.290 ;
    END
END AHHCINX2

MACRO AFHCONX2
    CLASS CORE ;
    FOREIGN AFHCONX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.460 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  20.090 0.650 20.330 4.300 ;
        RECT  19.900 0.650 20.090 1.550 ;
        RECT  19.900 2.380 20.090 4.300 ;
        RECT  19.250 2.380 19.900 3.780 ;
        END
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.540 1.990 13.940 2.390 ;
        RECT  13.350 3.480 13.750 3.880 ;
        RECT  12.150 2.080 13.540 2.320 ;
        RECT  12.160 3.510 13.350 3.750 ;
        RECT  11.760 3.430 12.160 3.830 ;
        RECT  11.250 1.920 12.150 2.320 ;
        RECT  11.670 3.510 11.760 3.830 ;
        RECT  11.430 3.510 11.670 3.750 ;
        RECT  11.330 3.510 11.430 3.780 ;
        RECT  11.110 3.500 11.330 3.780 ;
        RECT  11.110 2.080 11.250 2.320 ;
        RECT  10.870 2.080 11.110 3.780 ;
        RECT  10.670 2.380 10.870 3.780 ;
        END
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  18.280 1.990 18.340 2.390 ;
        RECT  18.020 1.990 18.280 2.650 ;
        RECT  17.940 1.990 18.020 2.390 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.040 1.840 9.560 2.240 ;
        RECT  8.780 1.830 9.040 2.240 ;
        RECT  8.160 1.840 8.780 2.240 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.330 2.070 1.870 2.660 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  19.580 4.640 20.460 5.440 ;
        RECT  19.180 4.180 19.580 5.440 ;
        RECT  17.440 4.640 19.180 5.440 ;
        RECT  17.040 4.480 17.440 5.440 ;
        RECT  9.320 4.640 17.040 5.440 ;
        RECT  8.920 4.480 9.320 5.440 ;
        RECT  1.350 4.640 8.920 5.440 ;
        RECT  0.950 4.480 1.350 5.440 ;
        RECT  0.000 4.640 0.950 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  19.580 -0.400 20.460 0.400 ;
        RECT  19.180 -0.400 19.580 0.780 ;
        RECT  17.300 -0.400 19.180 0.400 ;
        RECT  16.900 -0.400 17.300 0.560 ;
        RECT  9.320 -0.400 16.900 0.400 ;
        RECT  8.920 -0.400 9.320 0.560 ;
        RECT  1.350 -0.400 8.920 0.400 ;
        RECT  0.950 -0.400 1.350 0.560 ;
        RECT  0.000 -0.400 0.950 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  19.510 1.880 19.780 2.120 ;
        RECT  19.270 1.020 19.510 2.120 ;
        RECT  18.780 1.020 19.270 1.260 ;
        RECT  18.620 1.500 18.860 4.400 ;
        RECT  18.540 0.800 18.780 1.260 ;
        RECT  18.410 1.500 18.620 1.740 ;
        RECT  18.460 3.540 18.620 4.400 ;
        RECT  15.710 0.800 18.540 1.040 ;
        RECT  14.680 3.680 18.460 3.920 ;
        RECT  17.410 2.900 18.230 3.140 ;
        RECT  17.410 1.300 18.090 1.540 ;
        RECT  17.170 1.300 17.410 3.440 ;
        RECT  16.850 1.850 17.170 2.250 ;
        RECT  15.490 3.200 17.170 3.440 ;
        RECT  16.610 2.560 16.930 2.960 ;
        RECT  10.410 4.160 16.700 4.400 ;
        RECT  16.370 1.300 16.610 2.960 ;
        RECT  16.110 1.300 16.370 1.540 ;
        RECT  15.890 2.290 16.130 2.960 ;
        RECT  15.710 2.290 15.890 2.530 ;
        RECT  15.470 0.720 15.710 2.530 ;
        RECT  15.230 3.040 15.490 3.440 ;
        RECT  14.990 1.790 15.230 3.440 ;
        RECT  14.750 0.640 14.990 2.030 ;
        RECT  14.510 2.270 14.740 2.670 ;
        RECT  14.440 2.920 14.680 3.920 ;
        RECT  14.270 0.800 14.510 2.670 ;
        RECT  13.750 2.920 14.440 3.160 ;
        RECT  8.690 0.800 14.270 1.040 ;
        RECT  13.540 1.280 13.940 1.590 ;
        RECT  13.350 2.760 13.750 3.160 ;
        RECT  10.040 1.280 13.540 1.520 ;
        RECT  12.160 2.780 13.350 3.020 ;
        RECT  11.760 2.710 12.160 3.110 ;
        RECT  10.170 3.960 10.410 4.400 ;
        RECT  7.720 3.960 10.170 4.200 ;
        RECT  10.040 2.820 10.110 3.720 ;
        RECT  9.800 1.280 10.040 3.720 ;
        RECT  9.710 1.280 9.800 1.520 ;
        RECT  9.710 2.820 9.800 3.720 ;
        RECT  8.450 0.680 8.690 1.040 ;
        RECT  7.880 1.280 8.530 1.520 ;
        RECT  8.370 2.820 8.530 3.720 ;
        RECT  7.240 0.680 8.450 0.920 ;
        RECT  8.130 2.480 8.370 3.720 ;
        RECT  7.880 2.480 8.130 2.720 ;
        RECT  7.480 1.160 7.880 2.720 ;
        RECT  7.480 2.970 7.720 4.200 ;
        RECT  7.160 2.320 7.480 2.720 ;
        RECT  6.890 2.970 7.480 3.210 ;
        RECT  7.000 0.680 7.240 1.610 ;
        RECT  6.890 1.370 7.000 1.610 ;
        RECT  5.990 1.370 6.890 1.770 ;
        RECT  5.990 2.090 6.890 2.490 ;
        RECT  5.990 2.810 6.890 3.210 ;
        RECT  6.230 3.580 6.890 3.980 ;
        RECT  4.300 0.730 6.760 0.970 ;
        RECT  5.990 3.580 6.230 4.360 ;
        RECT  4.780 1.530 5.990 1.770 ;
        RECT  5.270 2.250 5.990 2.490 ;
        RECT  5.750 2.970 5.990 3.210 ;
        RECT  3.060 4.120 5.990 4.360 ;
        RECT  5.510 2.970 5.750 3.560 ;
        RECT  4.780 3.320 5.510 3.560 ;
        RECT  5.030 2.250 5.270 2.840 ;
        RECT  4.780 2.600 5.030 2.840 ;
        RECT  4.540 1.530 4.780 2.280 ;
        RECT  3.380 2.600 4.780 3.000 ;
        RECT  3.380 3.320 4.780 3.720 ;
        RECT  3.380 1.880 4.540 2.280 ;
        RECT  4.060 0.730 4.300 1.560 ;
        RECT  3.400 1.160 4.060 1.560 ;
        RECT  2.880 1.160 3.400 1.400 ;
        RECT  2.350 2.680 3.380 2.920 ;
        RECT  2.820 3.780 3.060 4.360 ;
        RECT  2.640 0.890 2.880 1.400 ;
        RECT  0.560 3.780 2.820 4.020 ;
        RECT  0.560 0.890 2.640 1.130 ;
        RECT  2.140 1.400 2.350 3.350 ;
        RECT  2.110 1.400 2.140 3.510 ;
        RECT  1.740 1.400 2.110 1.800 ;
        RECT  1.740 3.110 2.110 3.510 ;
        RECT  1.050 3.110 1.740 3.350 ;
        RECT  0.810 2.080 1.050 3.350 ;
        RECT  0.650 2.080 0.810 2.480 ;
        RECT  0.400 0.690 0.560 1.590 ;
        RECT  0.400 2.820 0.560 4.220 ;
        RECT  0.160 0.690 0.400 4.220 ;
    END
END AFHCONX2

MACRO AFHCINX2
    CLASS CORE ;
    FOREIGN AFHCINX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.980 1.250 18.210 3.490 ;
        RECT  17.810 0.690 17.980 3.490 ;
        RECT  17.580 0.690 17.810 1.650 ;
        RECT  17.800 3.090 17.810 3.490 ;
        RECT  17.370 3.090 17.800 4.340 ;
        RECT  17.270 3.500 17.370 4.340 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.570 1.280 11.730 1.680 ;
        RECT  11.330 1.280 11.570 2.060 ;
        RECT  11.130 1.820 11.330 2.060 ;
        RECT  10.890 1.820 11.130 3.760 ;
        RECT  10.670 1.820 10.890 2.660 ;
        END
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  13.060 2.180 13.070 2.580 ;
        RECT  12.680 2.180 13.060 2.660 ;
        RECT  12.670 2.180 12.680 2.580 ;
        END
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.710 4.060 7.720 4.340 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.010 2.950 1.120 3.210 ;
        RECT  0.770 2.160 1.010 3.210 ;
        RECT  0.650 2.170 0.770 2.570 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  16.340 4.640 18.480 5.440 ;
        RECT  15.940 4.480 16.340 5.440 ;
        RECT  13.030 4.640 15.940 5.440 ;
        RECT  12.630 4.480 13.030 5.440 ;
        RECT  9.670 4.640 12.630 5.440 ;
        RECT  9.270 4.480 9.670 5.440 ;
        RECT  1.280 4.640 9.270 5.440 ;
        RECT  0.880 3.570 1.280 5.440 ;
        RECT  0.000 4.640 0.880 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  17.190 -0.400 18.480 0.400 ;
        RECT  16.790 -0.400 17.190 0.560 ;
        RECT  13.260 -0.400 16.790 0.400 ;
        RECT  12.860 -0.400 13.260 0.560 ;
        RECT  9.270 -0.400 12.860 0.400 ;
        RECT  8.870 -0.400 9.270 0.560 ;
        RECT  1.350 -0.400 8.870 0.400 ;
        RECT  0.950 -0.400 1.350 0.560 ;
        RECT  0.000 -0.400 0.950 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  17.410 2.000 17.570 2.400 ;
        RECT  17.170 2.000 17.410 2.780 ;
        RECT  16.790 2.540 17.170 2.780 ;
        RECT  16.570 0.800 16.810 2.290 ;
        RECT  16.550 2.540 16.790 4.240 ;
        RECT  16.230 0.800 16.570 1.040 ;
        RECT  14.720 4.000 16.550 4.240 ;
        RECT  16.070 1.300 16.310 3.600 ;
        RECT  15.990 0.700 16.230 1.040 ;
        RECT  15.530 3.360 16.070 3.600 ;
        RECT  14.890 0.700 15.990 0.940 ;
        RECT  15.590 1.530 15.830 3.030 ;
        RECT  15.410 1.530 15.590 1.770 ;
        RECT  14.720 2.790 15.590 3.030 ;
        RECT  15.130 3.360 15.530 3.760 ;
        RECT  15.170 1.180 15.410 1.770 ;
        RECT  14.240 2.150 15.350 2.550 ;
        RECT  14.650 0.700 14.890 1.580 ;
        RECT  14.480 2.790 14.720 4.240 ;
        RECT  14.330 1.180 14.650 1.580 ;
        RECT  13.740 0.640 14.410 0.880 ;
        RECT  13.760 1.340 14.330 1.580 ;
        RECT  14.000 2.150 14.240 4.240 ;
        RECT  11.610 4.000 14.000 4.240 ;
        RECT  13.520 1.340 13.760 3.760 ;
        RECT  13.500 0.640 13.740 1.040 ;
        RECT  12.440 0.800 13.500 1.040 ;
        RECT  12.300 1.290 12.460 1.690 ;
        RECT  12.200 0.640 12.440 1.040 ;
        RECT  12.060 1.290 12.300 3.760 ;
        RECT  9.750 0.640 12.200 0.880 ;
        RECT  11.890 2.860 12.060 3.760 ;
        RECT  11.370 2.300 11.610 4.240 ;
        RECT  8.200 4.000 11.370 4.240 ;
        RECT  10.600 1.180 11.000 1.580 ;
        RECT  10.400 1.300 10.600 1.580 ;
        RECT  10.160 1.300 10.400 3.760 ;
        RECT  9.660 1.300 10.160 1.700 ;
        RECT  8.850 2.160 9.770 2.560 ;
        RECT  9.510 0.640 9.750 1.040 ;
        RECT  8.190 0.800 9.510 1.040 ;
        RECT  8.470 2.160 8.850 3.640 ;
        RECT  8.450 1.300 8.470 3.640 ;
        RECT  8.070 1.300 8.450 2.660 ;
        RECT  7.960 3.580 8.200 4.240 ;
        RECT  7.950 0.640 8.190 1.040 ;
        RECT  7.770 2.240 8.070 2.660 ;
        RECT  6.860 3.580 7.960 3.820 ;
        RECT  7.530 0.640 7.950 0.880 ;
        RECT  7.290 0.640 7.530 3.340 ;
        RECT  5.420 0.640 7.290 0.880 ;
        RECT  7.110 2.940 7.290 3.340 ;
        RECT  6.860 1.120 7.050 2.500 ;
        RECT  6.810 1.120 6.860 3.820 ;
        RECT  5.900 1.120 6.810 1.360 ;
        RECT  6.620 2.260 6.810 3.820 ;
        RECT  6.380 1.600 6.560 2.000 ;
        RECT  6.140 1.600 6.380 4.390 ;
        RECT  2.060 4.150 6.140 4.390 ;
        RECT  5.660 1.120 5.900 3.910 ;
        RECT  4.060 3.670 5.660 3.910 ;
        RECT  5.180 0.640 5.420 3.360 ;
        RECT  4.640 0.640 4.880 3.260 ;
        RECT  2.300 0.640 4.640 0.880 ;
        RECT  4.380 2.840 4.640 3.260 ;
        RECT  3.330 2.840 4.380 3.080 ;
        RECT  3.840 1.120 4.240 1.540 ;
        RECT  3.660 3.320 4.060 3.910 ;
        RECT  2.860 1.300 3.840 1.540 ;
        RECT  2.690 3.670 3.660 3.910 ;
        RECT  2.930 2.840 3.330 3.260 ;
        RECT  2.690 1.300 2.860 1.700 ;
        RECT  2.450 1.300 2.690 3.910 ;
        RECT  2.320 3.670 2.450 3.910 ;
        RECT  2.060 0.640 2.300 1.040 ;
        RECT  2.060 1.290 2.140 1.690 ;
        RECT  1.500 0.800 2.060 1.040 ;
        RECT  1.820 1.290 2.060 4.390 ;
        RECT  1.740 1.290 1.820 1.690 ;
        RECT  1.600 2.920 1.820 4.390 ;
        RECT  1.500 1.920 1.570 2.320 ;
        RECT  1.260 0.800 1.500 2.320 ;
        RECT  0.560 0.800 1.260 1.040 ;
        RECT  0.400 0.720 0.560 1.620 ;
        RECT  0.400 3.000 0.480 4.400 ;
        RECT  0.160 0.720 0.400 4.400 ;
    END
END AFHCINX2

MACRO CMPR42X2
    CLASS CORE ;
    FOREIGN CMPR42X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 26.400 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  25.840 2.660 25.880 3.640 ;
        RECT  25.880 2.380 25.950 3.640 ;
        RECT  25.840 0.970 25.950 1.370 ;
        RECT  25.950 0.970 26.190 3.640 ;
        RECT  26.190 2.380 26.220 3.640 ;
        RECT  26.220 2.640 26.240 3.640 ;
        RECT  26.190 0.970 26.240 1.370 ;
        END
    END S
    PIN ICO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.160 0.860 0.200 3.740 ;
        RECT  0.200 0.860 0.400 3.770 ;
        RECT  0.400 2.840 0.460 3.770 ;
        RECT  0.460 2.840 0.560 3.740 ;
        RECT  0.400 0.860 0.560 1.280 ;
        END
    END ICO
    PIN ICI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  22.550 1.380 22.990 2.180 ;
        END
    END ICI
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  14.540 2.560 14.700 2.800 ;
        RECT  14.700 2.080 14.940 2.800 ;
        RECT  14.940 2.080 16.700 2.320 ;
        RECT  16.700 1.830 16.960 2.320 ;
        RECT  16.960 2.080 17.500 2.320 ;
        END
    END D
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  20.120 3.140 20.510 3.380 ;
        RECT  20.110 1.180 20.510 1.420 ;
        RECT  20.510 1.180 20.750 3.380 ;
        RECT  20.750 2.950 20.920 3.210 ;
        END
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.240 4.000 3.650 4.400 ;
        RECT  3.650 4.000 6.830 4.240 ;
        RECT  6.830 4.000 7.070 4.400 ;
        RECT  7.070 4.160 8.860 4.400 ;
        RECT  8.860 4.000 9.100 4.400 ;
        RECT  9.100 4.000 10.760 4.240 ;
        RECT  10.760 4.000 11.020 4.330 ;
        RECT  11.020 4.000 14.140 4.240 ;
        RECT  14.140 4.000 14.380 4.400 ;
        RECT  14.380 4.160 17.200 4.400 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.970 2.340 3.440 2.580 ;
        RECT  3.440 2.340 3.500 2.640 ;
        RECT  3.500 2.340 3.760 2.650 ;
        RECT  3.760 2.340 3.830 2.640 ;
        RECT  3.830 2.340 5.070 2.580 ;
        RECT  5.070 2.340 5.140 2.660 ;
        RECT  5.140 2.340 5.380 3.760 ;
        RECT  5.380 3.520 6.370 3.760 ;
        RECT  6.370 2.720 6.610 3.760 ;
        RECT  6.610 2.720 7.420 2.960 ;
        RECT  7.420 2.520 7.660 2.960 ;
        RECT  7.660 2.520 8.480 2.760 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.330 1.800 1.570 2.500 ;
        RECT  1.570 1.800 1.780 2.090 ;
        RECT  1.780 1.800 3.910 2.040 ;
        RECT  3.910 1.760 4.310 2.040 ;
        RECT  4.310 1.760 6.350 2.000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.950 5.440 ;
        RECT  0.950 3.810 1.350 5.440 ;
        RECT  1.350 4.640 5.200 5.440 ;
        RECT  5.200 4.480 5.600 5.440 ;
        RECT  5.600 4.640 6.200 5.440 ;
        RECT  6.200 4.480 6.600 5.440 ;
        RECT  6.600 4.640 9.340 5.440 ;
        RECT  9.340 4.480 9.740 5.440 ;
        RECT  9.740 4.640 13.500 5.440 ;
        RECT  13.500 4.480 13.900 5.440 ;
        RECT  16.470 3.500 17.370 3.920 ;
        RECT  13.900 4.640 17.440 5.440 ;
        RECT  17.370 3.660 17.440 3.920 ;
        RECT  17.440 3.660 17.700 5.440 ;
        RECT  17.700 4.640 21.980 5.440 ;
        RECT  21.980 4.480 22.380 5.440 ;
        RECT  22.380 4.640 25.040 5.440 ;
        RECT  25.040 4.480 25.200 5.440 ;
        RECT  25.200 3.780 25.440 5.440 ;
        RECT  25.440 4.640 26.400 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.950 0.400 ;
        RECT  0.950 -0.400 1.350 0.560 ;
        RECT  1.350 -0.400 3.430 0.400 ;
        RECT  3.430 -0.400 3.830 0.560 ;
        RECT  3.830 -0.400 5.040 0.400 ;
        RECT  5.040 -0.400 5.440 0.560 ;
        RECT  5.440 -0.400 6.540 0.400 ;
        RECT  6.540 -0.400 6.940 0.560 ;
        RECT  6.940 -0.400 9.300 0.400 ;
        RECT  9.300 -0.400 9.700 0.560 ;
        RECT  9.700 -0.400 12.400 0.400 ;
        RECT  12.400 -0.400 12.800 0.560 ;
        RECT  12.800 -0.400 16.920 0.400 ;
        RECT  16.920 -0.400 17.320 0.560 ;
        RECT  17.320 -0.400 22.000 0.400 ;
        RECT  22.000 -0.400 22.400 0.560 ;
        RECT  22.400 -0.400 25.050 0.400 ;
        RECT  25.050 -0.400 25.450 0.560 ;
        RECT  25.450 -0.400 26.400 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  25.580 1.900 25.610 2.300 ;
        RECT  25.340 0.800 25.580 3.540 ;
        RECT  23.800 0.800 25.340 1.040 ;
        RECT  24.960 3.300 25.340 3.540 ;
        RECT  24.860 1.280 25.100 2.930 ;
        RECT  24.720 3.300 24.960 4.240 ;
        RECT  23.510 1.280 24.860 1.520 ;
        RECT  24.480 2.690 24.860 2.930 ;
        RECT  23.910 4.000 24.720 4.240 ;
        RECT  23.500 1.990 24.590 2.230 ;
        RECT  24.240 2.690 24.480 3.760 ;
        RECT  23.170 3.520 24.240 3.760 ;
        RECT  23.760 2.610 24.000 3.280 ;
        RECT  23.510 4.000 23.910 4.310 ;
        RECT  21.830 3.040 23.760 3.280 ;
        RECT  23.270 0.900 23.510 1.520 ;
        RECT  23.260 1.990 23.500 2.780 ;
        RECT  23.080 0.900 23.270 1.140 ;
        RECT  22.310 2.540 23.260 2.780 ;
        RECT  23.010 3.520 23.170 3.920 ;
        RECT  22.770 3.520 23.010 4.240 ;
        RECT  21.710 4.000 22.770 4.240 ;
        RECT  22.070 0.850 22.310 2.780 ;
        RECT  21.230 0.850 22.070 1.090 ;
        RECT  21.790 1.340 21.830 3.280 ;
        RECT  21.590 1.340 21.790 3.730 ;
        RECT  21.470 4.000 21.710 4.400 ;
        RECT  21.530 1.340 21.590 1.740 ;
        RECT  21.550 2.930 21.590 3.730 ;
        RECT  21.230 3.490 21.550 3.730 ;
        RECT  19.530 4.160 21.470 4.400 ;
        RECT  21.230 1.940 21.350 2.400 ;
        RECT  20.990 0.640 21.230 2.400 ;
        RECT  20.990 3.490 21.230 3.920 ;
        RECT  18.510 0.640 20.990 0.880 ;
        RECT  19.790 3.680 20.990 3.920 ;
        RECT  20.030 1.660 20.270 2.870 ;
        RECT  19.790 1.660 20.030 1.900 ;
        RECT  19.700 2.630 20.030 2.870 ;
        RECT  19.550 1.180 19.790 1.900 ;
        RECT  19.120 2.140 19.790 2.380 ;
        RECT  19.530 2.630 19.700 3.440 ;
        RECT  19.390 1.180 19.550 1.420 ;
        RECT  19.460 2.630 19.530 4.400 ;
        RECT  19.290 3.040 19.460 4.400 ;
        RECT  18.990 2.000 19.120 2.380 ;
        RECT  18.750 1.120 18.990 3.770 ;
        RECT  18.580 3.370 18.750 3.770 ;
        RECT  18.270 0.640 18.510 2.880 ;
        RECT  18.030 3.180 18.280 3.760 ;
        RECT  16.450 0.800 18.270 1.040 ;
        RECT  17.940 1.280 18.030 3.760 ;
        RECT  17.790 1.280 17.940 3.420 ;
        RECT  17.780 2.710 17.790 3.420 ;
        RECT  15.830 2.710 17.780 2.950 ;
        RECT  16.240 1.280 16.530 1.520 ;
        RECT  16.210 0.640 16.450 1.040 ;
        RECT  16.000 1.280 16.240 1.840 ;
        RECT  13.280 0.640 16.210 0.880 ;
        RECT  15.830 3.190 16.070 3.760 ;
        RECT  14.240 1.600 16.000 1.840 ;
        RECT  15.590 2.560 15.830 2.950 ;
        RECT  15.350 3.190 15.830 3.430 ;
        RECT  13.760 1.120 15.710 1.360 ;
        RECT  15.260 2.560 15.590 2.800 ;
        RECT  14.860 3.680 15.430 3.920 ;
        RECT  15.110 3.040 15.350 3.430 ;
        RECT  14.240 3.040 15.110 3.280 ;
        RECT  14.620 3.520 14.860 3.920 ;
        RECT  13.720 3.520 14.620 3.760 ;
        RECT  14.000 1.600 14.240 3.280 ;
        RECT  13.800 2.080 14.000 2.480 ;
        RECT  13.520 1.120 13.760 1.520 ;
        RECT  13.480 2.980 13.720 3.760 ;
        RECT  12.580 1.280 13.520 1.520 ;
        RECT  12.580 2.980 13.480 3.220 ;
        RECT  13.040 0.640 13.280 1.040 ;
        RECT  9.760 3.520 13.230 3.760 ;
        RECT  11.810 0.800 13.040 1.040 ;
        RECT  12.340 1.280 12.580 3.220 ;
        RECT  12.050 1.280 12.340 1.680 ;
        RECT  11.810 2.980 12.010 3.220 ;
        RECT  11.570 0.800 11.810 3.220 ;
        RECT  10.810 0.800 11.570 1.200 ;
        RECT  11.080 1.800 11.320 2.200 ;
        RECT  10.490 1.800 11.080 2.040 ;
        RECT  10.370 2.960 10.530 3.200 ;
        RECT  10.370 0.800 10.490 2.040 ;
        RECT  10.130 0.800 10.370 3.200 ;
        RECT  10.090 0.800 10.130 1.200 ;
        RECT  9.520 0.800 9.760 3.760 ;
        RECT  8.450 0.800 9.520 1.040 ;
        RECT  8.620 3.520 9.520 3.760 ;
        RECT  9.020 1.280 9.260 2.770 ;
        RECT  7.730 1.280 9.020 1.520 ;
        RECT  9.000 2.530 9.020 2.770 ;
        RECT  8.760 2.530 9.000 3.250 ;
        RECT  8.140 3.010 8.760 3.250 ;
        RECT  7.180 1.820 8.720 2.060 ;
        RECT  8.380 3.520 8.620 3.920 ;
        RECT  8.050 0.640 8.450 1.040 ;
        RECT  7.710 3.680 8.380 3.920 ;
        RECT  7.900 3.010 8.140 3.440 ;
        RECT  6.990 3.200 7.900 3.440 ;
        RECT  7.330 0.990 7.730 1.520 ;
        RECT  6.980 1.820 7.180 2.480 ;
        RECT  6.740 1.250 6.980 2.480 ;
        RECT  6.100 1.250 6.740 1.490 ;
        RECT  6.130 2.240 6.740 2.480 ;
        RECT  5.890 2.240 6.130 3.280 ;
        RECT  5.700 1.090 6.100 1.490 ;
        RECT  5.730 2.880 5.890 3.280 ;
        RECT  4.410 3.210 4.810 3.610 ;
        RECT  4.250 0.830 4.650 1.320 ;
        RECT  3.320 3.210 4.410 3.450 ;
        RECT  3.320 1.080 4.250 1.320 ;
        RECT  2.920 1.080 3.320 1.510 ;
        RECT  2.920 3.210 3.320 3.610 ;
        RECT  2.200 1.120 2.600 1.520 ;
        RECT  2.200 3.290 2.600 3.690 ;
        RECT  1.040 1.280 2.200 1.520 ;
        RECT  1.040 3.290 2.200 3.530 ;
        RECT  0.800 1.280 1.040 3.530 ;
        RECT  0.650 1.960 0.800 2.360 ;
    END
END CMPR42X2

MACRO CMPR42X1
    CLASS CORE ;
    FOREIGN CMPR42X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CMPR42X2 ;
    SIZE 23.100 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  22.540 2.390 22.700 3.390 ;
        RECT  22.540 1.170 22.700 1.570 ;
        RECT  22.700 1.170 22.940 3.390 ;
        END
    END S
    PIN ICO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.160 1.320 0.400 3.210 ;
        RECT  0.400 2.950 0.560 3.210 ;
        RECT  0.400 1.320 0.560 1.840 ;
        END
    END ICO
    PIN ICI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  19.240 2.290 19.690 3.080 ;
        END
    END ICI
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  12.840 1.660 13.080 2.100 ;
        RECT  13.080 1.820 13.940 2.100 ;
        RECT  13.940 1.820 14.180 2.340 ;
        END
    END D
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.050 2.880 17.130 3.280 ;
        RECT  16.970 1.180 17.130 1.580 ;
        RECT  17.130 1.180 17.370 3.280 ;
        RECT  17.370 1.830 17.620 2.090 ;
        END
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.850 4.160 5.700 4.400 ;
        RECT  5.700 4.000 6.150 4.400 ;
        RECT  6.150 4.000 8.180 4.240 ;
        RECT  8.180 4.000 8.420 4.400 ;
        RECT  8.420 4.160 9.510 4.400 ;
        RECT  9.510 4.000 9.750 4.400 ;
        RECT  9.750 4.000 12.650 4.240 ;
        RECT  12.650 3.500 12.750 4.240 ;
        RECT  12.750 3.500 13.090 4.300 ;
        RECT  13.090 4.060 13.400 4.300 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.060 2.270 3.500 2.510 ;
        RECT  3.500 2.270 3.760 2.650 ;
        RECT  3.760 2.270 4.190 2.610 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.340 1.780 1.780 2.400 ;
        RECT  1.780 1.780 4.550 2.020 ;
        RECT  4.550 1.780 4.790 2.480 ;
        RECT  4.790 2.080 4.870 2.480 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.920 5.440 ;
        RECT  0.920 4.480 1.320 5.440 ;
        RECT  1.320 4.640 2.500 5.440 ;
        RECT  2.500 4.480 3.370 5.440 ;
        RECT  3.370 3.680 3.610 5.440 ;
        RECT  3.610 3.680 4.850 3.920 ;
        RECT  4.850 3.410 5.250 3.920 ;
        RECT  3.610 4.640 7.420 5.440 ;
        RECT  7.420 4.480 7.820 5.440 ;
        RECT  7.820 4.640 10.700 5.440 ;
        RECT  10.700 4.480 11.100 5.440 ;
        RECT  11.100 4.640 13.640 5.440 ;
        RECT  13.640 3.170 14.040 5.440 ;
        RECT  14.040 4.640 17.560 5.440 ;
        RECT  17.560 4.480 17.960 5.440 ;
        RECT  17.960 4.640 18.890 5.440 ;
        RECT  18.890 3.810 19.290 5.440 ;
        RECT  19.290 4.640 22.300 5.440 ;
        RECT  22.300 4.480 22.700 5.440 ;
        RECT  22.700 4.640 23.100 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.750 0.400 ;
        RECT  0.750 -0.400 1.150 0.560 ;
        RECT  1.150 -0.400 3.590 0.400 ;
        RECT  3.590 -0.400 3.990 0.560 ;
        RECT  3.990 -0.400 4.840 0.400 ;
        RECT  4.840 -0.400 5.240 1.040 ;
        RECT  5.240 -0.400 7.600 0.400 ;
        RECT  7.600 -0.400 8.000 0.560 ;
        RECT  8.000 -0.400 10.550 0.400 ;
        RECT  10.550 -0.400 10.950 0.560 ;
        RECT  10.950 -0.400 13.820 0.400 ;
        RECT  13.820 -0.400 14.220 0.560 ;
        RECT  14.220 -0.400 18.260 0.400 ;
        RECT  18.260 -0.400 18.660 0.560 ;
        RECT  18.660 -0.400 21.810 0.400 ;
        RECT  21.810 -0.400 22.050 1.260 ;
        RECT  22.050 -0.400 22.440 0.560 ;
        RECT  22.440 -0.400 23.100 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  22.120 2.400 22.240 2.800 ;
        RECT  21.880 1.500 22.120 4.080 ;
        RECT  21.550 1.500 21.880 1.740 ;
        RECT  20.810 3.840 21.880 4.080 ;
        RECT  21.360 1.980 21.600 3.570 ;
        RECT  21.310 0.740 21.550 1.740 ;
        RECT  21.100 1.980 21.360 2.380 ;
        RECT  20.050 3.330 21.360 3.570 ;
        RECT  20.120 0.740 21.310 0.980 ;
        RECT  20.970 1.980 21.100 2.220 ;
        RECT  20.210 2.850 21.060 3.090 ;
        RECT  20.730 1.220 20.970 2.220 ;
        RECT  20.410 3.810 20.810 4.080 ;
        RECT  19.660 1.220 20.730 1.460 ;
        RECT  19.970 1.700 20.210 3.090 ;
        RECT  19.650 3.330 20.050 3.960 ;
        RECT  18.830 1.700 19.970 1.940 ;
        RECT  19.420 0.640 19.660 1.460 ;
        RECT  18.560 3.330 19.650 3.570 ;
        RECT  19.260 0.640 19.420 1.040 ;
        RECT  18.590 1.400 18.830 3.090 ;
        RECT  18.500 1.400 18.590 1.800 ;
        RECT  18.420 2.800 18.590 3.090 ;
        RECT  18.320 3.330 18.560 4.240 ;
        RECT  17.950 2.850 18.420 3.090 ;
        RECT  18.190 2.000 18.350 2.400 ;
        RECT  16.270 4.000 18.320 4.240 ;
        RECT  17.950 1.230 18.190 2.400 ;
        RECT  17.710 0.640 17.950 1.470 ;
        RECT  17.710 2.850 17.950 3.760 ;
        RECT  15.200 0.640 17.710 0.880 ;
        RECT  16.750 3.520 17.710 3.760 ;
        RECT  16.510 3.360 16.750 3.760 ;
        RECT  16.480 1.210 16.720 3.000 ;
        RECT  16.220 1.210 16.480 1.610 ;
        RECT  16.270 2.760 16.480 3.000 ;
        RECT  16.030 2.760 16.270 4.240 ;
        RECT  16.000 2.110 16.240 2.510 ;
        RECT  15.870 3.470 16.030 3.870 ;
        RECT  15.680 2.110 16.000 2.350 ;
        RECT  15.550 1.210 15.680 3.220 ;
        RECT  15.440 1.210 15.550 3.840 ;
        RECT  15.310 2.980 15.440 3.840 ;
        RECT  15.150 3.440 15.310 3.840 ;
        RECT  14.960 0.640 15.200 2.720 ;
        RECT  14.750 0.640 14.960 1.040 ;
        RECT  14.900 2.320 14.960 2.720 ;
        RECT  14.660 3.520 14.830 3.760 ;
        RECT  13.580 0.800 14.750 1.040 ;
        RECT  14.660 1.280 14.720 1.680 ;
        RECT  14.420 1.280 14.660 3.760 ;
        RECT  13.700 2.580 14.420 2.820 ;
        RECT  13.460 2.420 13.700 2.820 ;
        RECT  13.340 0.640 13.580 1.040 ;
        RECT  12.180 2.420 13.460 2.660 ;
        RECT  11.510 0.640 13.340 0.880 ;
        RECT  12.600 1.120 13.090 1.360 ;
        RECT  12.670 2.960 13.070 3.260 ;
        RECT  11.930 2.960 12.670 3.200 ;
        RECT  12.360 1.120 12.600 2.180 ;
        RECT  11.930 1.940 12.360 2.180 ;
        RECT  11.950 3.440 12.350 3.760 ;
        RECT  11.880 1.120 12.120 1.700 ;
        RECT  10.640 3.520 11.950 3.760 ;
        RECT  11.690 1.940 11.930 3.200 ;
        RECT  11.410 1.460 11.880 1.700 ;
        RECT  11.400 2.310 11.690 2.550 ;
        RECT  11.270 0.640 11.510 1.220 ;
        RECT  11.170 1.460 11.410 1.840 ;
        RECT  11.000 2.230 11.400 2.630 ;
        RECT  10.590 0.980 11.270 1.220 ;
        RECT  10.640 1.600 11.170 1.840 ;
        RECT  10.400 1.600 10.640 3.760 ;
        RECT  10.350 0.980 10.590 1.360 ;
        RECT  9.920 1.600 10.400 1.840 ;
        RECT  10.230 2.160 10.400 2.560 ;
        RECT  10.160 3.200 10.400 3.600 ;
        RECT  9.680 1.120 10.350 1.360 ;
        RECT  8.780 0.640 9.940 0.880 ;
        RECT  9.680 3.200 9.840 3.600 ;
        RECT  9.440 1.120 9.680 3.600 ;
        RECT  9.100 1.300 9.440 1.700 ;
        RECT  8.720 3.520 9.120 3.920 ;
        RECT  8.540 0.640 8.780 3.200 ;
        RECT  7.910 3.520 8.720 3.760 ;
        RECT  8.380 1.300 8.540 1.700 ;
        RECT  8.210 2.960 8.540 3.200 ;
        RECT  8.140 2.060 8.270 2.460 ;
        RECT  7.910 1.090 8.140 2.720 ;
        RECT  7.900 1.090 7.910 3.760 ;
        RECT  6.750 1.090 7.900 1.330 ;
        RECT  7.670 2.480 7.900 3.760 ;
        RECT  6.710 3.520 7.670 3.760 ;
        RECT  6.960 2.000 7.660 2.240 ;
        RECT  6.720 1.670 6.960 3.070 ;
        RECT  6.350 0.930 6.750 1.330 ;
        RECT  6.030 1.670 6.720 1.910 ;
        RECT  5.910 2.830 6.720 3.070 ;
        RECT  6.310 3.320 6.710 3.760 ;
        RECT  6.080 2.170 6.480 2.570 ;
        RECT  5.350 2.170 6.080 2.560 ;
        RECT  5.790 0.900 6.030 1.910 ;
        RECT  5.670 2.830 5.910 3.470 ;
        RECT  5.630 0.900 5.790 1.300 ;
        RECT  5.110 1.280 5.350 3.170 ;
        RECT  4.600 1.280 5.110 1.520 ;
        RECT  4.380 2.930 5.110 3.170 ;
        RECT  3.980 1.120 4.600 1.520 ;
        RECT  3.980 2.930 4.380 3.370 ;
        RECT  3.350 1.300 3.590 1.540 ;
        RECT  3.120 2.950 3.410 3.190 ;
        RECT  3.110 0.640 3.350 1.540 ;
        RECT  2.880 2.950 3.120 4.210 ;
        RECT  1.610 0.640 3.110 0.880 ;
        RECT  2.110 3.970 2.880 4.210 ;
        RECT  2.470 1.120 2.870 1.540 ;
        RECT  2.370 2.860 2.610 3.260 ;
        RECT  1.090 1.120 2.470 1.360 ;
        RECT  1.090 2.860 2.370 3.100 ;
        RECT  1.710 3.970 2.110 4.370 ;
        RECT  0.850 0.810 1.090 3.100 ;
        RECT  0.510 0.810 0.850 1.050 ;
        RECT  0.270 0.640 0.510 1.050 ;
    END
END CMPR42X1

MACRO BMXX1
    CLASS CORE ;
    FOREIGN BMXX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN X2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.380 2.260 9.840 2.820 ;
        RECT  9.840 2.420 9.870 2.820 ;
        END
    END X2
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.730 2.180 7.140 2.670 ;
        END
    END S
    PIN PP
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.980 3.220 12.060 3.690 ;
        RECT  12.060 1.230 12.300 3.690 ;
        RECT  12.300 2.950 12.340 3.690 ;
        RECT  12.340 3.200 12.380 3.690 ;
        END
    END PP
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.030 1.840 6.140 2.410 ;
        RECT  6.140 1.830 6.400 2.410 ;
        RECT  6.400 1.840 6.430 2.410 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.640 2.060 0.770 2.460 ;
        RECT  0.770 1.820 1.040 2.460 ;
        RECT  1.040 1.820 1.110 2.090 ;
        RECT  1.110 1.830 1.120 2.090 ;
        END
    END M0
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.470 2.170 1.520 2.570 ;
        RECT  1.520 2.170 1.780 2.650 ;
        RECT  1.780 2.170 1.870 2.570 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.000 5.440 ;
        RECT  1.000 3.860 1.400 5.440 ;
        RECT  1.400 4.640 6.490 5.440 ;
        RECT  6.490 4.480 6.890 5.440 ;
        RECT  6.890 4.640 8.590 5.440 ;
        RECT  8.590 4.480 9.490 5.440 ;
        RECT  9.490 4.640 11.560 5.440 ;
        RECT  11.560 4.480 11.960 5.440 ;
        RECT  11.960 4.640 12.540 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.020 0.400 ;
        RECT  1.020 -0.400 1.420 1.500 ;
        RECT  1.420 -0.400 6.270 0.400 ;
        RECT  6.270 -0.400 7.670 0.560 ;
        RECT  7.670 -0.400 11.710 0.400 ;
        RECT  11.710 -0.400 12.110 0.560 ;
        RECT  12.110 -0.400 12.540 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  11.530 1.210 11.750 3.050 ;
        RECT  11.510 1.210 11.530 4.240 ;
        RECT  11.470 1.210 11.510 1.450 ;
        RECT  11.310 2.810 11.510 4.240 ;
        RECT  11.230 0.640 11.470 1.450 ;
        RECT  11.290 2.810 11.310 4.400 ;
        RECT  11.070 4.000 11.290 4.400 ;
        RECT  10.380 2.160 11.270 2.560 ;
        RECT  9.720 0.640 11.230 0.880 ;
        RECT  9.900 4.160 11.070 4.400 ;
        RECT  10.830 3.250 11.020 3.650 ;
        RECT  10.750 1.120 10.990 1.900 ;
        RECT  10.590 3.250 10.830 3.890 ;
        RECT  8.630 1.120 10.750 1.360 ;
        RECT  8.630 3.650 10.590 3.890 ;
        RECT  10.350 1.600 10.380 2.560 ;
        RECT  10.110 1.600 10.350 3.380 ;
        RECT  9.950 1.600 10.110 1.840 ;
        RECT  9.900 3.140 10.110 3.380 ;
        RECT  9.110 1.600 9.630 1.840 ;
        RECT  9.110 3.100 9.580 3.340 ;
        RECT  8.150 0.640 9.330 0.880 ;
        RECT  8.870 1.600 9.110 3.340 ;
        RECT  8.390 1.120 8.630 1.630 ;
        RECT  8.390 3.260 8.630 3.890 ;
        RECT  8.120 1.390 8.390 1.630 ;
        RECT  8.120 3.260 8.390 3.500 ;
        RECT  7.910 0.640 8.150 1.040 ;
        RECT  5.950 4.000 8.150 4.240 ;
        RECT  7.880 1.390 8.120 3.500 ;
        RECT  5.990 0.800 7.910 1.040 ;
        RECT  7.480 1.500 7.630 3.410 ;
        RECT  7.400 1.420 7.480 3.570 ;
        RECT  7.390 1.420 7.400 3.760 ;
        RECT  7.080 1.420 7.390 1.820 ;
        RECT  7.080 3.170 7.390 3.760 ;
        RECT  5.470 3.520 7.080 3.760 ;
        RECT  5.790 2.720 6.100 3.120 ;
        RECT  5.790 1.330 6.030 1.570 ;
        RECT  5.750 0.780 5.990 1.040 ;
        RECT  5.710 4.000 5.950 4.400 ;
        RECT  5.700 1.330 5.790 3.120 ;
        RECT  4.510 0.780 5.750 1.020 ;
        RECT  3.010 4.160 5.710 4.400 ;
        RECT  5.550 1.330 5.700 3.040 ;
        RECT  5.230 2.020 5.550 2.420 ;
        RECT  5.230 3.520 5.470 3.920 ;
        RECT  4.990 1.260 5.310 1.500 ;
        RECT  4.990 2.700 5.300 3.100 ;
        RECT  3.550 3.680 5.230 3.920 ;
        RECT  4.750 1.260 4.990 3.440 ;
        RECT  4.030 3.200 4.750 3.440 ;
        RECT  4.270 0.780 4.510 2.960 ;
        RECT  3.790 0.700 4.030 3.440 ;
        RECT  2.350 0.700 3.790 0.940 ;
        RECT  3.310 1.180 3.550 3.920 ;
        RECT  2.830 2.900 3.010 4.400 ;
        RECT  2.770 1.180 2.830 4.400 ;
        RECT  2.590 1.180 2.770 3.140 ;
        RECT  2.120 3.380 2.520 3.860 ;
        RECT  2.110 0.700 2.350 3.140 ;
        RECT  0.560 3.380 2.120 3.620 ;
        RECT  1.790 1.180 2.110 1.580 ;
        RECT  1.790 2.900 2.110 3.140 ;
        RECT  0.400 2.720 0.560 3.620 ;
        RECT  0.400 1.420 0.480 1.820 ;
        RECT  0.320 1.420 0.400 3.620 ;
        RECT  0.160 1.420 0.320 3.120 ;
    END
END BMXX1

MACRO BENCX4
    CLASS CORE ;
    FOREIGN BENCX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 48.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN X2
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  28.850 2.900 32.130 3.140 ;
        RECT  32.130 2.900 32.450 3.220 ;
        RECT  28.180 1.280 32.450 1.520 ;
        RECT  32.450 1.280 32.890 3.220 ;
        RECT  32.890 2.900 33.210 3.220 ;
        RECT  32.890 1.280 33.380 1.520 ;
        RECT  33.210 2.900 34.080 3.140 ;
        END
    END X2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  42.720 0.810 42.800 1.770 ;
        RECT  42.690 2.800 43.090 3.760 ;
        RECT  43.090 2.800 43.110 3.220 ;
        RECT  42.800 0.810 43.120 1.830 ;
        RECT  43.110 2.800 44.010 3.040 ;
        RECT  44.010 2.800 44.130 3.220 ;
        RECT  43.120 1.590 44.160 1.830 ;
        RECT  44.130 2.800 44.530 3.760 ;
        RECT  44.160 0.810 44.560 1.830 ;
        RECT  44.530 2.800 45.330 3.040 ;
        RECT  45.330 2.800 45.570 3.220 ;
        RECT  44.560 1.590 45.600 1.830 ;
        RECT  45.570 2.800 45.970 3.760 ;
        RECT  45.600 0.810 46.000 1.830 ;
        RECT  45.970 2.800 46.650 3.040 ;
        RECT  46.650 2.800 46.970 3.220 ;
        RECT  46.000 1.590 46.970 1.830 ;
        RECT  46.970 1.540 47.010 3.220 ;
        RECT  47.010 1.540 47.040 3.760 ;
        RECT  47.040 0.810 47.410 3.760 ;
        RECT  47.410 0.810 47.440 3.140 ;
        END
    END S
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  16.480 4.000 16.700 4.240 ;
        RECT  16.700 4.000 16.960 4.330 ;
        RECT  16.960 4.000 21.810 4.240 ;
        RECT  21.810 4.000 22.050 4.390 ;
        RECT  22.050 4.150 25.890 4.390 ;
        RECT  25.890 4.000 26.130 4.390 ;
        RECT  26.130 4.000 35.690 4.240 ;
        END
    END M2
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  10.010 2.490 10.250 3.530 ;
        RECT  10.250 3.200 10.450 3.530 ;
        RECT  10.450 3.290 11.800 3.530 ;
        RECT  11.800 2.580 12.200 3.530 ;
        RECT  12.200 3.200 12.430 3.530 ;
        RECT  12.430 3.290 13.770 3.530 ;
        RECT  13.770 3.290 14.010 3.750 ;
        RECT  14.010 3.510 14.310 3.750 ;
        RECT  14.310 3.510 14.410 3.780 ;
        RECT  14.410 3.500 15.020 3.780 ;
        RECT  15.020 3.500 15.260 4.250 ;
        RECT  15.260 3.500 15.270 4.170 ;
        RECT  15.270 3.500 15.290 3.780 ;
        RECT  15.290 3.520 21.870 3.760 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  10.650 2.520 10.670 2.760 ;
        RECT  10.670 2.060 11.050 2.760 ;
        RECT  11.050 2.060 11.110 2.660 ;
        RECT  11.110 2.060 14.290 2.300 ;
        RECT  14.290 0.800 14.530 2.300 ;
        RECT  14.530 0.800 15.660 1.040 ;
        RECT  15.660 0.650 15.900 1.040 ;
        RECT  15.900 0.650 16.620 0.890 ;
        RECT  16.620 0.650 16.860 2.260 ;
        RECT  16.860 2.020 18.260 2.260 ;
        END
    END M0
    PIN A
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.880 0.850 1.070 1.970 ;
        RECT  1.070 0.850 1.280 4.190 ;
        RECT  1.280 1.570 1.470 4.190 ;
        RECT  1.470 1.570 1.870 3.220 ;
        RECT  1.870 2.730 2.190 3.220 ;
        RECT  1.870 1.570 2.330 1.810 ;
        RECT  2.190 2.730 2.430 2.970 ;
        RECT  2.430 2.730 2.520 3.220 ;
        RECT  2.330 0.850 2.730 1.810 ;
        RECT  2.520 2.730 2.920 4.190 ;
        RECT  2.920 2.730 3.750 2.970 ;
        RECT  2.730 1.570 3.790 1.810 ;
        RECT  3.750 2.730 3.990 3.220 ;
        RECT  3.790 0.850 4.190 1.810 ;
        RECT  3.990 2.730 4.390 4.190 ;
        RECT  4.190 1.570 5.240 1.810 ;
        RECT  4.390 2.730 5.440 2.970 ;
        RECT  5.240 0.850 5.640 1.810 ;
        RECT  5.440 2.730 5.840 4.190 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.350 5.440 ;
        RECT  0.350 2.730 0.750 5.440 ;
        RECT  0.750 4.640 1.790 5.440 ;
        RECT  1.790 3.530 2.190 5.440 ;
        RECT  2.190 4.640 3.270 5.440 ;
        RECT  3.270 3.490 3.670 5.440 ;
        RECT  3.670 4.640 4.720 5.440 ;
        RECT  4.720 3.530 5.120 5.440 ;
        RECT  5.120 4.640 6.160 5.440 ;
        RECT  6.160 3.530 6.560 5.440 ;
        RECT  6.560 4.640 7.610 5.440 ;
        RECT  7.610 3.530 8.010 5.440 ;
        RECT  8.010 4.640 9.630 5.440 ;
        RECT  9.630 4.480 10.030 5.440 ;
        RECT  10.030 4.640 12.130 5.440 ;
        RECT  12.130 4.480 12.530 5.440 ;
        RECT  12.530 4.640 14.380 5.440 ;
        RECT  14.380 4.060 14.780 5.440 ;
        RECT  14.780 4.640 15.840 5.440 ;
        RECT  15.840 4.060 16.240 5.440 ;
        RECT  16.240 4.640 17.570 5.440 ;
        RECT  17.570 4.480 17.970 5.440 ;
        RECT  17.970 4.640 19.220 5.440 ;
        RECT  19.220 4.480 19.620 5.440 ;
        RECT  19.620 4.640 20.750 5.440 ;
        RECT  20.750 4.480 21.150 5.440 ;
        RECT  21.150 4.640 26.480 5.440 ;
        RECT  26.480 4.480 26.880 5.440 ;
        RECT  26.880 4.640 28.060 5.440 ;
        RECT  28.060 4.480 28.460 5.440 ;
        RECT  28.460 4.640 29.650 5.440 ;
        RECT  29.650 4.480 30.050 5.440 ;
        RECT  30.050 4.640 31.260 5.440 ;
        RECT  31.260 4.480 31.660 5.440 ;
        RECT  31.660 4.640 32.890 5.440 ;
        RECT  32.890 4.480 33.290 5.440 ;
        RECT  33.290 4.640 34.500 5.440 ;
        RECT  34.500 4.480 34.900 5.440 ;
        RECT  34.900 4.640 36.420 5.440 ;
        RECT  36.420 4.480 36.820 5.440 ;
        RECT  36.820 4.640 39.010 5.440 ;
        RECT  39.010 4.480 39.410 5.440 ;
        RECT  39.410 4.640 40.390 5.440 ;
        RECT  40.390 3.520 40.790 5.440 ;
        RECT  40.790 4.640 41.970 5.440 ;
        RECT  41.970 3.540 42.370 5.440 ;
        RECT  42.370 4.640 43.410 5.440 ;
        RECT  43.410 3.490 43.810 5.440 ;
        RECT  43.810 4.640 44.850 5.440 ;
        RECT  44.850 3.540 45.250 5.440 ;
        RECT  45.250 4.640 46.290 5.440 ;
        RECT  46.290 3.490 46.690 5.440 ;
        RECT  46.690 4.640 47.730 5.440 ;
        RECT  47.730 3.540 48.130 5.440 ;
        RECT  48.130 4.640 48.840 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 1.610 ;
        RECT  0.560 -0.400 1.610 0.400 ;
        RECT  1.610 -0.400 2.010 1.060 ;
        RECT  2.010 -0.400 3.060 0.400 ;
        RECT  3.060 -0.400 3.460 1.060 ;
        RECT  3.460 -0.400 4.510 0.400 ;
        RECT  4.510 -0.400 4.910 1.060 ;
        RECT  4.910 -0.400 5.960 0.400 ;
        RECT  5.960 -0.400 6.360 1.190 ;
        RECT  6.360 -0.400 7.400 0.400 ;
        RECT  7.400 -0.400 7.800 1.190 ;
        RECT  7.800 -0.400 8.660 0.400 ;
        RECT  8.660 -0.400 9.060 1.030 ;
        RECT  9.060 -0.400 10.170 0.400 ;
        RECT  10.170 -0.400 10.570 0.560 ;
        RECT  10.570 -0.400 11.770 0.400 ;
        RECT  11.770 -0.400 12.170 0.560 ;
        RECT  12.170 -0.400 15.010 0.400 ;
        RECT  15.010 -0.400 15.410 0.560 ;
        RECT  15.410 -0.400 17.740 0.400 ;
        RECT  17.740 -0.400 18.140 1.000 ;
        RECT  18.140 -0.400 19.250 0.400 ;
        RECT  19.250 -0.400 19.650 0.560 ;
        RECT  19.650 -0.400 25.920 0.400 ;
        RECT  25.920 -0.400 26.320 0.560 ;
        RECT  26.320 -0.400 27.360 0.400 ;
        RECT  27.360 -0.400 27.760 0.560 ;
        RECT  27.760 -0.400 28.990 0.400 ;
        RECT  28.990 -0.400 29.390 0.560 ;
        RECT  29.390 -0.400 30.590 0.400 ;
        RECT  30.590 -0.400 30.990 0.560 ;
        RECT  30.990 -0.400 32.190 0.400 ;
        RECT  32.190 -0.400 32.590 0.560 ;
        RECT  32.590 -0.400 33.790 0.400 ;
        RECT  33.790 -0.400 34.190 0.560 ;
        RECT  34.190 -0.400 36.300 0.400 ;
        RECT  36.300 -0.400 36.700 0.560 ;
        RECT  36.700 -0.400 37.850 0.400 ;
        RECT  37.850 -0.400 38.250 0.560 ;
        RECT  38.250 -0.400 39.360 0.400 ;
        RECT  39.360 -0.400 39.600 0.980 ;
        RECT  39.600 -0.400 40.520 0.400 ;
        RECT  40.520 -0.400 40.920 1.210 ;
        RECT  40.920 -0.400 42.000 0.400 ;
        RECT  42.000 -0.400 42.400 1.210 ;
        RECT  42.400 -0.400 43.440 0.400 ;
        RECT  43.440 -0.400 43.840 1.300 ;
        RECT  43.840 -0.400 44.880 0.400 ;
        RECT  44.880 -0.400 45.280 1.290 ;
        RECT  45.280 -0.400 46.320 0.400 ;
        RECT  46.320 -0.400 46.720 1.300 ;
        RECT  46.720 -0.400 47.760 0.400 ;
        RECT  47.760 -0.400 48.160 1.530 ;
        RECT  48.160 -0.400 48.840 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  42.350 2.270 46.410 2.510 ;
        RECT  42.110 1.450 42.350 3.070 ;
        RECT  39.790 1.450 42.110 1.690 ;
        RECT  41.510 2.830 42.110 3.070 ;
        RECT  40.280 2.090 41.740 2.490 ;
        RECT  41.110 2.830 41.510 3.790 ;
        RECT  40.070 2.830 41.110 3.070 ;
        RECT  39.380 2.100 40.280 2.490 ;
        RECT  39.670 2.830 40.070 3.790 ;
        RECT  39.140 1.660 39.380 3.660 ;
        RECT  36.310 1.660 39.140 1.900 ;
        RECT  35.620 3.420 39.140 3.660 ;
        RECT  36.830 1.180 38.960 1.420 ;
        RECT  38.660 2.570 38.900 3.120 ;
        RECT  37.120 2.880 38.660 3.120 ;
        RECT  38.230 2.390 38.300 2.630 ;
        RECT  37.900 2.160 38.230 2.630 ;
        RECT  33.860 2.160 37.900 2.400 ;
        RECT  36.720 2.660 37.120 3.120 ;
        RECT  36.590 0.880 36.830 1.420 ;
        RECT  34.850 2.880 36.720 3.120 ;
        RECT  35.060 0.880 36.590 1.120 ;
        RECT  36.070 1.380 36.310 1.900 ;
        RECT  34.650 1.380 36.070 1.620 ;
        RECT  34.610 2.880 34.850 3.740 ;
        RECT  34.410 1.220 34.650 1.620 ;
        RECT  26.210 3.500 34.610 3.740 ;
        RECT  33.620 0.800 33.860 2.400 ;
        RECT  25.540 0.800 33.620 1.040 ;
        RECT  27.670 2.080 32.080 2.320 ;
        RECT  27.430 1.360 27.670 3.040 ;
        RECT  25.130 1.360 27.430 1.600 ;
        RECT  27.270 2.710 27.430 3.040 ;
        RECT  25.660 2.710 27.270 2.950 ;
        RECT  26.070 2.170 27.140 2.410 ;
        RECT  25.970 3.190 26.210 3.740 ;
        RECT  25.830 1.890 26.070 2.410 ;
        RECT  25.330 3.190 25.970 3.430 ;
        RECT  24.740 1.890 25.830 2.130 ;
        RECT  22.540 3.670 25.550 3.910 ;
        RECT  25.300 0.640 25.540 1.040 ;
        RECT  25.090 2.400 25.330 3.430 ;
        RECT  23.860 0.640 25.300 0.880 ;
        RECT  24.740 1.140 24.810 1.380 ;
        RECT  24.500 1.140 24.740 3.430 ;
        RECT  24.410 1.140 24.500 1.380 ;
        RECT  23.140 3.190 24.500 3.430 ;
        RECT  23.860 2.710 24.020 2.950 ;
        RECT  23.620 0.640 23.860 2.950 ;
        RECT  21.010 0.640 23.620 0.880 ;
        RECT  23.140 1.120 23.370 1.360 ;
        RECT  22.900 1.120 23.140 3.430 ;
        RECT  21.390 1.120 22.900 1.360 ;
        RECT  22.540 1.600 22.580 1.840 ;
        RECT  22.300 1.600 22.540 3.910 ;
        RECT  21.060 1.600 22.300 1.840 ;
        RECT  22.180 3.040 22.300 3.540 ;
        RECT  19.950 3.040 22.180 3.280 ;
        RECT  19.520 2.560 22.060 2.800 ;
        RECT  20.820 1.380 21.060 1.840 ;
        RECT  20.770 0.640 21.010 1.040 ;
        RECT  20.060 1.380 20.820 1.620 ;
        RECT  19.660 0.800 20.770 1.040 ;
        RECT  19.660 1.940 19.970 2.180 ;
        RECT  19.420 0.800 19.660 2.180 ;
        RECT  19.280 2.560 19.520 3.280 ;
        RECT  18.860 1.320 19.420 1.560 ;
        RECT  16.380 3.040 19.280 3.280 ;
        RECT  18.760 1.160 18.860 1.560 ;
        RECT  18.520 1.160 18.760 2.800 ;
        RECT  18.460 1.160 18.520 1.560 ;
        RECT  16.810 2.560 18.520 2.800 ;
        RECT  17.340 1.320 18.460 1.560 ;
        RECT  17.100 1.160 17.340 1.560 ;
        RECT  16.140 1.180 16.380 3.280 ;
        RECT  15.260 2.700 16.140 3.100 ;
        RECT  14.770 1.280 15.010 3.010 ;
        RECT  13.120 2.770 14.770 3.010 ;
        RECT  13.810 0.950 14.050 1.520 ;
        RECT  12.690 0.950 13.810 1.190 ;
        RECT  13.330 1.430 13.410 1.670 ;
        RECT  9.720 3.780 13.390 4.020 ;
        RECT  13.010 1.430 13.330 1.790 ;
        RECT  12.880 2.660 13.120 3.010 ;
        RECT  9.720 1.550 13.010 1.790 ;
        RECT  12.690 2.660 12.880 2.900 ;
        RECT  12.370 0.950 12.690 1.290 ;
        RECT  9.380 1.050 12.370 1.290 ;
        RECT  9.480 1.550 9.720 4.020 ;
        RECT  6.660 2.070 9.480 2.470 ;
        RECT  8.330 3.050 8.730 4.010 ;
        RECT  6.330 1.430 8.530 1.670 ;
        RECT  7.290 3.050 8.330 3.290 ;
        RECT  6.890 3.050 7.290 4.010 ;
        RECT  6.330 3.050 6.890 3.290 ;
        RECT  6.090 1.430 6.330 3.290 ;
        RECT  2.110 2.150 6.090 2.390 ;
    END
END BENCX4

MACRO XOR3X4
    CLASS CORE ;
    FOREIGN XOR3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.120 2.900 17.270 4.300 ;
        RECT  17.270 2.900 17.370 4.340 ;
        RECT  17.120 0.790 17.370 1.690 ;
        RECT  17.370 0.790 17.520 4.340 ;
        RECT  17.520 1.440 17.610 4.340 ;
        RECT  17.610 2.940 17.710 4.340 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  15.380 4.070 15.690 4.330 ;
        RECT  15.690 3.980 15.830 4.330 ;
        RECT  15.830 3.970 16.090 4.330 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.440 1.830 9.450 2.090 ;
        RECT  9.450 1.740 9.680 2.090 ;
        RECT  9.680 1.740 10.080 3.160 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.820 0.710 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.620 0.560 5.440 ;
        RECT  0.560 4.640 4.010 5.440 ;
        RECT  4.010 4.200 4.410 5.440 ;
        RECT  4.410 4.640 5.650 5.440 ;
        RECT  5.650 4.200 6.050 5.440 ;
        RECT  6.050 4.640 7.890 5.440 ;
        RECT  7.890 4.480 8.290 5.440 ;
        RECT  8.290 4.640 16.330 5.440 ;
        RECT  16.330 4.480 16.350 5.440 ;
        RECT  16.350 3.890 16.750 5.440 ;
        RECT  16.750 4.640 17.950 5.440 ;
        RECT  17.950 3.080 18.190 5.440 ;
        RECT  18.190 4.640 18.480 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 1.490 ;
        RECT  0.560 -0.400 4.300 0.400 ;
        RECT  4.300 -0.400 4.700 0.560 ;
        RECT  4.700 -0.400 5.880 0.400 ;
        RECT  5.880 -0.400 6.280 0.560 ;
        RECT  6.280 -0.400 16.400 0.400 ;
        RECT  16.400 -0.400 16.800 1.560 ;
        RECT  16.800 -0.400 17.850 0.400 ;
        RECT  17.850 -0.400 18.250 1.560 ;
        RECT  18.250 -0.400 18.480 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  17.050 2.100 17.130 2.500 ;
        RECT  16.880 2.100 17.050 2.660 ;
        RECT  16.730 2.100 16.880 3.600 ;
        RECT  16.640 2.420 16.730 3.600 ;
        RECT  15.720 3.360 16.640 3.600 ;
        RECT  15.560 1.420 15.960 3.120 ;
        RECT  15.480 3.360 15.720 3.700 ;
        RECT  15.030 2.180 15.560 2.580 ;
        RECT  14.520 3.460 15.480 3.700 ;
        RECT  14.840 2.820 15.240 3.220 ;
        RECT  14.760 1.120 14.890 1.520 ;
        RECT  14.760 2.820 14.840 3.060 ;
        RECT  14.730 1.120 14.760 3.060 ;
        RECT  14.520 0.640 14.730 3.060 ;
        RECT  14.490 0.640 14.520 1.520 ;
        RECT  14.280 3.300 14.520 3.700 ;
        RECT  11.920 0.640 14.490 0.880 ;
        RECT  14.170 1.790 14.280 3.700 ;
        RECT  14.120 1.120 14.170 3.700 ;
        RECT  14.040 1.120 14.120 3.550 ;
        RECT  13.930 1.120 14.040 2.030 ;
        RECT  13.770 1.120 13.930 1.520 ;
        RECT  13.410 3.040 13.800 3.940 ;
        RECT  12.740 1.120 13.770 1.360 ;
        RECT  13.170 1.600 13.410 4.400 ;
        RECT  12.980 1.600 13.170 1.840 ;
        RECT  8.810 4.160 13.170 4.400 ;
        RECT  12.740 3.040 12.920 3.920 ;
        RECT  12.500 1.120 12.740 3.920 ;
        RECT  12.190 1.120 12.500 1.520 ;
        RECT  11.920 3.040 12.080 3.920 ;
        RECT  11.680 0.640 11.920 3.920 ;
        RECT  11.470 0.710 11.680 1.820 ;
        RECT  10.560 0.710 11.470 0.950 ;
        RECT  11.070 3.240 11.360 3.640 ;
        RECT  10.830 1.410 11.070 3.920 ;
        RECT  9.290 3.680 10.830 3.920 ;
        RECT  10.320 0.710 10.560 3.440 ;
        RECT  10.030 0.980 10.320 1.500 ;
        RECT  8.610 1.260 10.030 1.500 ;
        RECT  8.130 0.780 9.500 1.020 ;
        RECT  9.200 2.480 9.440 3.130 ;
        RECT  9.050 3.520 9.290 3.920 ;
        RECT  8.610 2.480 9.200 2.720 ;
        RECT  7.650 3.520 9.050 3.760 ;
        RECT  8.570 4.000 8.810 4.400 ;
        RECT  8.130 2.960 8.800 3.200 ;
        RECT  8.370 1.260 8.610 2.720 ;
        RECT  7.650 4.000 8.570 4.240 ;
        RECT  7.890 0.780 8.130 3.200 ;
        RECT  5.970 0.800 7.890 1.040 ;
        RECT  7.410 1.280 7.650 3.760 ;
        RECT  7.410 4.000 7.650 4.400 ;
        RECT  6.450 1.280 7.410 1.520 ;
        RECT  6.530 4.160 7.410 4.400 ;
        RECT  7.150 3.680 7.170 3.920 ;
        RECT  6.770 1.760 7.150 3.920 ;
        RECT  6.750 1.760 6.770 3.480 ;
        RECT  3.190 3.240 6.750 3.480 ;
        RECT  6.290 3.720 6.530 4.400 ;
        RECT  6.210 1.280 6.450 3.000 ;
        RECT  3.670 3.720 6.290 3.960 ;
        RECT  5.110 2.760 6.210 3.000 ;
        RECT  5.750 0.800 5.970 2.410 ;
        RECT  5.730 0.800 5.750 2.490 ;
        RECT  4.060 0.900 5.730 1.140 ;
        RECT  5.350 2.090 5.730 2.490 ;
        RECT  5.110 1.380 5.490 1.840 ;
        RECT  5.090 1.380 5.110 3.000 ;
        RECT  4.870 1.600 5.090 3.000 ;
        RECT  2.710 1.600 4.870 1.840 ;
        RECT  3.820 0.640 4.060 1.140 ;
        RECT  1.200 0.640 3.820 0.880 ;
        RECT  3.430 3.720 3.670 4.180 ;
        RECT  1.680 1.120 3.580 1.360 ;
        RECT  1.680 3.940 3.430 4.180 ;
        RECT  2.950 3.240 3.190 3.700 ;
        RECT  2.160 3.460 2.950 3.700 ;
        RECT  2.470 1.600 2.710 3.220 ;
        RECT  2.390 1.600 2.470 1.840 ;
        RECT  1.920 2.180 2.160 3.700 ;
        RECT  1.440 1.120 1.680 4.180 ;
        RECT  0.960 0.640 1.200 4.220 ;
        RECT  0.950 0.640 0.960 1.420 ;
    END
END XOR3X4

MACRO XOR3X2
    CLASS CORE ;
    FOREIGN XOR3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ XOR3X4 ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.320 2.720 11.430 3.620 ;
        RECT  11.430 2.640 11.480 3.620 ;
        RECT  11.320 0.790 11.480 1.690 ;
        RECT  11.480 0.790 11.720 3.620 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  10.030 3.370 10.380 3.970 ;
        RECT  10.380 3.370 10.470 3.680 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.380 1.630 6.620 2.060 ;
        RECT  6.620 1.820 6.800 2.060 ;
        RECT  6.800 1.820 6.960 2.090 ;
        RECT  6.960 1.820 7.200 3.140 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.820 0.460 2.650 ;
        RECT  0.460 1.820 0.700 2.510 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.530 0.560 5.440 ;
        RECT  0.560 4.640 3.280 5.440 ;
        RECT  3.280 4.200 3.680 5.440 ;
        RECT  3.680 4.640 10.610 5.440 ;
        RECT  10.610 4.480 10.690 5.440 ;
        RECT  10.690 3.900 10.930 5.440 ;
        RECT  10.930 4.480 11.010 5.440 ;
        RECT  11.010 4.640 11.880 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 1.490 ;
        RECT  0.560 -0.400 3.410 0.400 ;
        RECT  3.410 -0.400 3.810 0.840 ;
        RECT  3.810 -0.400 10.530 0.400 ;
        RECT  10.530 -0.400 10.930 0.610 ;
        RECT  10.930 -0.400 11.880 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  11.020 1.950 11.200 2.350 ;
        RECT  10.780 0.850 11.020 2.350 ;
        RECT  10.140 0.850 10.780 1.090 ;
        RECT  10.180 1.470 10.300 1.710 ;
        RECT  10.180 2.720 10.300 3.120 ;
        RECT  9.900 1.470 10.180 3.120 ;
        RECT  9.900 0.680 10.140 1.090 ;
        RECT  8.820 0.680 9.900 0.920 ;
        RECT  9.780 1.930 9.900 2.330 ;
        RECT  9.540 3.680 9.770 4.400 ;
        RECT  9.520 1.260 9.540 4.400 ;
        RECT  9.300 1.180 9.520 4.400 ;
        RECT  9.120 1.180 9.300 1.580 ;
        RECT  4.160 4.160 9.300 4.400 ;
        RECT  8.820 2.890 9.060 3.790 ;
        RECT  8.660 0.680 8.820 3.790 ;
        RECT  8.580 0.680 8.660 3.140 ;
        RECT  8.400 0.930 8.580 1.330 ;
        RECT  8.160 3.270 8.340 3.670 ;
        RECT  7.920 0.860 8.160 3.670 ;
        RECT  7.640 0.860 7.920 1.100 ;
        RECT  7.620 1.340 7.680 3.820 ;
        RECT  7.400 0.640 7.640 1.100 ;
        RECT  7.440 1.340 7.620 3.900 ;
        RECT  7.100 1.340 7.440 1.580 ;
        RECT  7.220 3.500 7.440 3.900 ;
        RECT  6.300 0.640 7.400 0.880 ;
        RECT  5.180 3.500 7.220 3.740 ;
        RECT  6.860 1.120 7.100 1.580 ;
        RECT  6.620 1.120 6.860 1.360 ;
        RECT  6.560 2.780 6.720 3.180 ;
        RECT  6.320 2.340 6.560 3.180 ;
        RECT  6.140 2.340 6.320 2.580 ;
        RECT  6.140 0.640 6.300 1.320 ;
        RECT  6.060 0.640 6.140 2.580 ;
        RECT  5.900 0.920 6.060 2.580 ;
        RECT  5.660 2.820 6.000 3.220 ;
        RECT  5.600 1.050 5.660 3.220 ;
        RECT  5.520 1.050 5.600 3.110 ;
        RECT  5.420 0.920 5.520 3.110 ;
        RECT  5.120 0.920 5.420 1.320 ;
        RECT  4.940 1.560 5.180 3.740 ;
        RECT  3.170 1.080 5.120 1.320 ;
        RECT  3.730 1.560 4.940 1.800 ;
        RECT  4.640 2.040 4.700 2.280 ;
        RECT  4.400 2.040 4.640 3.680 ;
        RECT  4.300 2.040 4.400 2.900 ;
        RECT  2.180 3.240 4.400 3.480 ;
        RECT  4.210 2.500 4.300 2.900 ;
        RECT  3.920 3.720 4.160 4.400 ;
        RECT  1.700 3.720 3.920 3.960 ;
        RECT  3.490 1.560 3.730 3.000 ;
        RECT  2.690 2.760 3.490 3.000 ;
        RECT  2.930 0.700 3.170 2.310 ;
        RECT  1.200 0.700 2.930 0.940 ;
        RECT  2.450 1.180 2.690 3.000 ;
        RECT  2.420 2.760 2.450 3.000 ;
        RECT  1.940 2.080 2.180 3.480 ;
        RECT  1.890 1.180 2.050 1.580 ;
        RECT  1.700 1.180 1.890 1.840 ;
        RECT  1.650 1.180 1.700 3.960 ;
        RECT  1.460 1.600 1.650 3.960 ;
        RECT  0.960 0.700 1.200 4.280 ;
    END
END XOR3X2

MACRO XNOR3X4
    CLASS CORE ;
    FOREIGN XNOR3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.120 2.900 17.270 4.300 ;
        RECT  17.270 2.900 17.370 4.340 ;
        RECT  17.120 0.790 17.370 1.690 ;
        RECT  17.370 0.790 17.520 4.340 ;
        RECT  17.520 1.440 17.610 4.340 ;
        RECT  17.610 2.940 17.710 4.340 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  16.040 1.830 16.400 2.440 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.440 1.830 9.450 2.090 ;
        RECT  9.450 1.740 9.680 2.090 ;
        RECT  9.680 1.740 10.080 3.160 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.820 0.710 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.620 0.560 5.440 ;
        RECT  0.560 4.640 4.010 5.440 ;
        RECT  4.010 4.200 4.410 5.440 ;
        RECT  4.410 4.640 5.650 5.440 ;
        RECT  5.650 4.200 6.050 5.440 ;
        RECT  6.050 4.640 7.890 5.440 ;
        RECT  7.890 4.480 8.290 5.440 ;
        RECT  8.290 4.640 16.330 5.440 ;
        RECT  16.330 4.480 16.350 5.440 ;
        RECT  16.350 3.890 16.750 5.440 ;
        RECT  16.750 4.640 17.950 5.440 ;
        RECT  17.950 3.080 18.190 5.440 ;
        RECT  18.190 4.640 18.480 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 1.490 ;
        RECT  0.560 -0.400 4.300 0.400 ;
        RECT  4.300 -0.400 4.700 0.560 ;
        RECT  4.700 -0.400 5.880 0.400 ;
        RECT  5.880 -0.400 6.280 0.560 ;
        RECT  6.280 -0.400 16.400 0.400 ;
        RECT  16.400 -0.400 16.800 1.560 ;
        RECT  16.800 -0.400 17.850 0.400 ;
        RECT  17.850 -0.400 18.250 1.560 ;
        RECT  18.250 -0.400 18.480 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  17.050 2.100 17.130 2.500 ;
        RECT  16.880 2.100 17.050 2.660 ;
        RECT  16.730 2.100 16.880 3.600 ;
        RECT  16.640 2.420 16.730 3.600 ;
        RECT  15.720 3.360 16.640 3.600 ;
        RECT  15.710 1.180 16.010 1.580 ;
        RECT  15.800 2.720 15.960 3.120 ;
        RECT  15.710 2.340 15.800 3.120 ;
        RECT  15.480 3.360 15.720 4.200 ;
        RECT  15.610 1.180 15.710 3.120 ;
        RECT  15.560 1.340 15.610 3.120 ;
        RECT  15.470 1.340 15.560 2.580 ;
        RECT  14.520 3.960 15.480 4.200 ;
        RECT  15.070 1.760 15.470 2.160 ;
        RECT  15.080 2.820 15.240 3.720 ;
        RECT  14.840 2.470 15.080 3.720 ;
        RECT  14.830 1.120 14.890 1.520 ;
        RECT  14.830 2.470 14.840 2.710 ;
        RECT  14.730 1.120 14.830 2.710 ;
        RECT  14.590 0.640 14.730 2.710 ;
        RECT  14.490 0.640 14.590 1.520 ;
        RECT  14.350 3.050 14.520 4.200 ;
        RECT  11.920 0.640 14.490 0.880 ;
        RECT  14.280 1.790 14.350 4.200 ;
        RECT  14.170 1.790 14.280 3.950 ;
        RECT  14.110 1.120 14.170 3.950 ;
        RECT  13.930 1.120 14.110 2.030 ;
        RECT  13.770 1.120 13.930 1.520 ;
        RECT  13.410 3.040 13.800 3.940 ;
        RECT  12.740 1.120 13.770 1.360 ;
        RECT  13.170 1.600 13.410 4.400 ;
        RECT  12.980 1.600 13.170 1.840 ;
        RECT  8.810 4.160 13.170 4.400 ;
        RECT  12.740 3.040 12.920 3.920 ;
        RECT  12.500 1.120 12.740 3.920 ;
        RECT  12.190 1.120 12.500 1.520 ;
        RECT  11.920 3.040 12.080 3.920 ;
        RECT  11.680 0.640 11.920 3.920 ;
        RECT  11.470 0.710 11.680 1.820 ;
        RECT  10.560 0.710 11.470 0.950 ;
        RECT  11.070 3.240 11.360 3.640 ;
        RECT  10.830 1.410 11.070 3.920 ;
        RECT  9.290 3.680 10.830 3.920 ;
        RECT  10.320 0.710 10.560 3.440 ;
        RECT  10.030 0.980 10.320 1.500 ;
        RECT  8.610 1.260 10.030 1.500 ;
        RECT  8.130 0.780 9.500 1.020 ;
        RECT  9.200 2.480 9.440 3.130 ;
        RECT  9.050 3.520 9.290 3.920 ;
        RECT  8.610 2.480 9.200 2.720 ;
        RECT  7.650 3.520 9.050 3.760 ;
        RECT  8.570 4.000 8.810 4.400 ;
        RECT  8.130 2.960 8.800 3.200 ;
        RECT  8.370 1.260 8.610 2.720 ;
        RECT  7.650 4.000 8.570 4.240 ;
        RECT  7.890 0.780 8.130 3.200 ;
        RECT  5.970 0.800 7.890 1.040 ;
        RECT  7.410 1.280 7.650 3.760 ;
        RECT  7.410 4.000 7.650 4.400 ;
        RECT  6.450 1.280 7.410 1.520 ;
        RECT  6.530 4.160 7.410 4.400 ;
        RECT  7.150 3.680 7.170 3.920 ;
        RECT  6.770 1.760 7.150 3.920 ;
        RECT  6.750 1.760 6.770 3.480 ;
        RECT  3.190 3.240 6.750 3.480 ;
        RECT  6.290 3.720 6.530 4.400 ;
        RECT  6.210 1.280 6.450 3.000 ;
        RECT  3.670 3.720 6.290 3.960 ;
        RECT  5.110 2.760 6.210 3.000 ;
        RECT  5.750 0.800 5.970 2.410 ;
        RECT  5.730 0.800 5.750 2.490 ;
        RECT  4.060 0.900 5.730 1.140 ;
        RECT  5.350 2.090 5.730 2.490 ;
        RECT  5.110 1.380 5.490 1.840 ;
        RECT  5.090 1.380 5.110 3.000 ;
        RECT  4.870 1.600 5.090 3.000 ;
        RECT  2.710 1.600 4.870 1.840 ;
        RECT  3.820 0.640 4.060 1.140 ;
        RECT  1.200 0.640 3.820 0.880 ;
        RECT  3.430 3.720 3.670 4.180 ;
        RECT  1.680 1.120 3.580 1.360 ;
        RECT  1.680 3.940 3.430 4.180 ;
        RECT  2.950 3.240 3.190 3.700 ;
        RECT  2.160 3.460 2.950 3.700 ;
        RECT  2.470 1.600 2.710 3.220 ;
        RECT  2.390 1.600 2.470 1.840 ;
        RECT  1.920 2.180 2.160 3.700 ;
        RECT  1.440 1.120 1.680 4.180 ;
        RECT  0.960 0.640 1.200 4.220 ;
        RECT  0.950 0.640 0.960 1.420 ;
    END
END XNOR3X4

MACRO XNOR3X2
    CLASS CORE ;
    FOREIGN XNOR3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ XNOR3X4 ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.320 2.720 11.480 3.620 ;
        RECT  11.320 0.790 11.480 1.690 ;
        RECT  11.480 0.790 11.720 3.620 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  10.030 3.380 10.380 3.980 ;
        RECT  10.380 3.380 10.470 3.690 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.380 1.630 6.620 2.060 ;
        RECT  6.620 1.820 6.800 2.060 ;
        RECT  6.800 1.820 6.960 2.090 ;
        RECT  6.960 1.820 7.200 3.140 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.820 0.460 2.650 ;
        RECT  0.460 1.820 0.550 2.510 ;
        RECT  0.550 2.110 0.700 2.510 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.530 0.560 5.440 ;
        RECT  0.560 4.640 3.280 5.440 ;
        RECT  3.280 4.200 3.680 5.440 ;
        RECT  3.680 4.640 10.610 5.440 ;
        RECT  10.610 4.480 10.690 5.440 ;
        RECT  10.690 3.890 10.930 5.440 ;
        RECT  10.930 4.480 11.010 5.440 ;
        RECT  11.010 4.640 11.880 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 1.490 ;
        RECT  0.560 -0.400 3.410 0.400 ;
        RECT  3.410 -0.400 3.810 0.840 ;
        RECT  3.810 -0.400 10.530 0.400 ;
        RECT  10.530 -0.400 10.930 0.610 ;
        RECT  10.930 -0.400 11.880 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  11.020 1.950 11.200 2.350 ;
        RECT  10.780 0.930 11.020 2.350 ;
        RECT  10.140 0.930 10.780 1.170 ;
        RECT  10.180 1.410 10.300 1.810 ;
        RECT  10.180 2.720 10.300 3.120 ;
        RECT  9.900 1.410 10.180 3.120 ;
        RECT  9.900 0.680 10.140 1.170 ;
        RECT  8.820 0.680 9.900 0.920 ;
        RECT  9.880 1.410 9.900 2.580 ;
        RECT  9.780 2.180 9.880 2.580 ;
        RECT  9.540 3.680 9.770 4.400 ;
        RECT  9.520 1.260 9.540 4.400 ;
        RECT  9.300 1.180 9.520 4.400 ;
        RECT  9.120 1.180 9.300 1.580 ;
        RECT  4.160 4.160 9.300 4.400 ;
        RECT  8.820 2.890 9.060 3.790 ;
        RECT  8.660 0.680 8.820 3.790 ;
        RECT  8.580 0.680 8.660 3.140 ;
        RECT  8.400 0.680 8.580 1.580 ;
        RECT  8.160 3.270 8.340 3.670 ;
        RECT  7.920 0.860 8.160 3.670 ;
        RECT  7.640 0.860 7.920 1.100 ;
        RECT  7.620 1.340 7.680 3.820 ;
        RECT  7.400 0.640 7.640 1.100 ;
        RECT  7.440 1.340 7.620 3.900 ;
        RECT  7.100 1.340 7.440 1.580 ;
        RECT  7.220 3.500 7.440 3.900 ;
        RECT  6.300 0.640 7.400 0.880 ;
        RECT  5.180 3.500 7.220 3.740 ;
        RECT  6.860 1.120 7.100 1.580 ;
        RECT  6.620 1.120 6.860 1.360 ;
        RECT  6.560 2.780 6.720 3.180 ;
        RECT  6.320 2.340 6.560 3.180 ;
        RECT  6.140 2.340 6.320 2.580 ;
        RECT  6.140 0.640 6.300 1.320 ;
        RECT  6.060 0.640 6.140 2.580 ;
        RECT  5.900 0.920 6.060 2.580 ;
        RECT  5.660 2.820 6.000 3.220 ;
        RECT  5.600 1.050 5.660 3.220 ;
        RECT  5.520 1.050 5.600 3.110 ;
        RECT  5.420 0.920 5.520 3.110 ;
        RECT  5.120 0.920 5.420 1.320 ;
        RECT  4.940 1.560 5.180 3.740 ;
        RECT  3.170 1.080 5.120 1.320 ;
        RECT  3.730 1.560 4.940 1.800 ;
        RECT  4.640 2.040 4.700 2.280 ;
        RECT  4.400 2.040 4.640 3.680 ;
        RECT  4.300 2.040 4.400 2.900 ;
        RECT  2.180 3.240 4.400 3.480 ;
        RECT  4.210 2.500 4.300 2.900 ;
        RECT  3.920 3.720 4.160 4.400 ;
        RECT  1.700 3.720 3.920 3.960 ;
        RECT  3.490 1.560 3.730 3.000 ;
        RECT  2.690 2.760 3.490 3.000 ;
        RECT  2.930 0.700 3.170 2.310 ;
        RECT  1.200 0.700 2.930 0.940 ;
        RECT  2.450 1.180 2.690 3.000 ;
        RECT  2.420 2.760 2.450 3.000 ;
        RECT  1.940 2.080 2.180 3.480 ;
        RECT  1.890 1.180 2.050 1.580 ;
        RECT  1.700 1.180 1.890 1.840 ;
        RECT  1.650 1.180 1.700 3.960 ;
        RECT  1.460 1.600 1.650 3.960 ;
        RECT  0.960 0.700 1.200 4.280 ;
    END
END XNOR3X2

MACRO AFHCONX4
    CLASS CORE ;
    FOREIGN AFHCONX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AFHCONX2 ;
    SIZE 22.440 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.920 0.650 21.990 2.620 ;
        RECT  21.750 0.650 21.920 4.220 ;
        RECT  21.590 0.650 21.750 1.550 ;
        RECT  21.520 2.380 21.750 4.220 ;
        RECT  21.230 2.380 21.520 3.780 ;
        END
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.800 2.040 14.700 2.440 ;
        RECT  13.800 3.480 14.700 3.880 ;
        RECT  12.600 2.120 13.800 2.360 ;
        RECT  13.650 3.480 13.800 3.800 ;
        RECT  12.750 3.560 13.650 3.800 ;
        RECT  11.110 3.360 12.750 3.800 ;
        RECT  11.110 1.920 12.600 2.360 ;
        RECT  10.870 1.920 11.110 3.800 ;
        RECT  10.670 2.380 10.870 3.800 ;
        END
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  18.940 1.990 19.770 2.390 ;
        RECT  18.680 1.990 18.940 2.650 ;
        RECT  18.370 1.990 18.680 2.390 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.040 1.840 9.560 2.240 ;
        RECT  8.780 1.830 9.040 2.240 ;
        RECT  8.160 1.840 8.780 2.240 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.330 2.070 1.870 2.660 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  21.200 4.640 22.440 5.440 ;
        RECT  20.800 4.180 21.200 5.440 ;
        RECT  19.750 4.640 20.800 5.440 ;
        RECT  19.350 4.180 19.750 5.440 ;
        RECT  18.240 4.640 19.350 5.440 ;
        RECT  17.840 4.480 18.240 5.440 ;
        RECT  9.330 4.640 17.840 5.440 ;
        RECT  8.930 4.480 9.330 5.440 ;
        RECT  1.350 4.640 8.930 5.440 ;
        RECT  0.950 4.480 1.350 5.440 ;
        RECT  0.000 4.640 0.950 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  21.200 -0.400 22.440 0.400 ;
        RECT  20.800 -0.400 21.200 0.560 ;
        RECT  19.620 -0.400 20.800 0.400 ;
        RECT  19.220 -0.400 19.620 0.560 ;
        RECT  17.970 -0.400 19.220 0.400 ;
        RECT  17.570 -0.400 17.970 0.560 ;
        RECT  9.330 -0.400 17.570 0.400 ;
        RECT  8.930 -0.400 9.330 0.560 ;
        RECT  1.350 -0.400 8.930 0.400 ;
        RECT  0.950 -0.400 1.350 0.560 ;
        RECT  0.000 -0.400 0.950 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  20.890 1.880 21.500 2.120 ;
        RECT  20.650 0.800 20.890 2.120 ;
        RECT  16.380 0.800 20.650 1.040 ;
        RECT  20.410 3.250 20.470 4.150 ;
        RECT  20.070 1.300 20.410 4.150 ;
        RECT  20.010 1.300 20.070 3.900 ;
        RECT  15.350 3.580 20.010 3.820 ;
        RECT  18.080 2.940 19.030 3.340 ;
        RECT  18.080 1.300 18.830 1.540 ;
        RECT  17.840 1.300 18.080 3.340 ;
        RECT  17.600 1.850 17.840 2.250 ;
        RECT  16.160 3.100 17.840 3.340 ;
        RECT  17.360 2.620 17.600 2.860 ;
        RECT  10.410 4.160 17.370 4.400 ;
        RECT  17.120 1.300 17.360 2.860 ;
        RECT  16.780 1.300 17.120 1.540 ;
        RECT  16.660 2.620 16.880 2.860 ;
        RECT  16.420 1.780 16.660 2.860 ;
        RECT  16.380 1.780 16.420 2.020 ;
        RECT  16.140 0.720 16.380 2.020 ;
        RECT  15.900 2.940 16.160 3.340 ;
        RECT  15.660 1.790 15.900 3.340 ;
        RECT  15.420 0.640 15.660 2.030 ;
        RECT  15.180 2.270 15.410 2.670 ;
        RECT  15.110 2.920 15.350 3.820 ;
        RECT  14.940 0.800 15.180 2.670 ;
        RECT  14.700 2.920 15.110 3.160 ;
        RECT  13.850 0.800 14.940 1.040 ;
        RECT  13.800 1.280 14.700 1.720 ;
        RECT  13.800 2.760 14.700 3.160 ;
        RECT  13.450 0.790 13.850 1.040 ;
        RECT  10.040 1.280 13.800 1.520 ;
        RECT  12.780 2.840 13.800 3.080 ;
        RECT  8.690 0.800 13.450 1.040 ;
        RECT  11.380 2.640 12.780 3.080 ;
        RECT  10.170 3.960 10.410 4.400 ;
        RECT  7.720 3.960 10.170 4.200 ;
        RECT  10.040 2.820 10.120 3.720 ;
        RECT  9.800 1.280 10.040 3.720 ;
        RECT  9.720 1.280 9.800 1.520 ;
        RECT  9.720 2.820 9.800 3.720 ;
        RECT  8.450 0.680 8.690 1.040 ;
        RECT  7.880 1.280 8.540 1.520 ;
        RECT  8.380 2.820 8.540 3.720 ;
        RECT  7.240 0.680 8.450 0.920 ;
        RECT  8.140 2.480 8.380 3.720 ;
        RECT  7.880 2.480 8.140 2.720 ;
        RECT  7.480 1.160 7.880 2.720 ;
        RECT  7.480 2.970 7.720 4.200 ;
        RECT  7.160 2.320 7.480 2.720 ;
        RECT  6.890 2.970 7.480 3.210 ;
        RECT  7.000 0.680 7.240 1.610 ;
        RECT  6.890 1.370 7.000 1.610 ;
        RECT  5.990 1.370 6.890 1.770 ;
        RECT  5.990 2.090 6.890 2.490 ;
        RECT  5.990 2.810 6.890 3.210 ;
        RECT  6.230 3.580 6.890 3.980 ;
        RECT  4.300 0.730 6.760 0.970 ;
        RECT  5.990 3.580 6.230 4.360 ;
        RECT  4.780 1.530 5.990 1.770 ;
        RECT  5.270 2.250 5.990 2.490 ;
        RECT  5.750 2.970 5.990 3.210 ;
        RECT  3.060 4.120 5.990 4.360 ;
        RECT  5.510 2.970 5.750 3.560 ;
        RECT  4.780 3.320 5.510 3.560 ;
        RECT  5.030 2.250 5.270 2.840 ;
        RECT  4.780 2.600 5.030 2.840 ;
        RECT  4.540 1.530 4.780 2.280 ;
        RECT  3.380 2.600 4.780 3.000 ;
        RECT  3.380 3.320 4.780 3.720 ;
        RECT  3.380 1.880 4.540 2.280 ;
        RECT  4.060 0.730 4.300 1.560 ;
        RECT  3.400 1.160 4.060 1.560 ;
        RECT  2.880 1.160 3.400 1.400 ;
        RECT  2.350 2.680 3.380 2.920 ;
        RECT  2.820 3.780 3.060 4.360 ;
        RECT  2.640 0.890 2.880 1.400 ;
        RECT  0.560 3.780 2.820 4.020 ;
        RECT  0.560 0.890 2.640 1.130 ;
        RECT  2.140 1.400 2.350 3.350 ;
        RECT  2.110 1.400 2.140 3.510 ;
        RECT  1.740 1.400 2.110 1.800 ;
        RECT  1.740 3.110 2.110 3.510 ;
        RECT  1.050 3.110 1.740 3.350 ;
        RECT  0.810 2.080 1.050 3.350 ;
        RECT  0.650 2.080 0.810 2.480 ;
        RECT  0.400 0.690 0.560 1.590 ;
        RECT  0.400 2.820 0.560 4.220 ;
        RECT  0.160 0.690 0.400 4.220 ;
    END
END AFHCONX4

MACRO AFHCINX4
    CLASS CORE ;
    FOREIGN AFHCINX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AFHCINX2 ;
    SIZE 23.100 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.970 1.600 14.410 3.280 ;
        RECT  13.950 2.880 13.970 3.280 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.810 2.280 22.330 3.900 ;
        RECT  21.770 1.130 21.810 3.900 ;
        RECT  21.570 1.130 21.770 2.620 ;
        RECT  20.730 3.660 21.770 3.900 ;
        RECT  21.410 1.130 21.570 1.530 ;
        RECT  20.330 2.940 20.730 3.900 ;
        RECT  19.980 2.940 20.330 3.180 ;
        RECT  19.740 1.760 19.980 3.180 ;
        RECT  19.580 1.760 19.740 2.000 ;
        END
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  17.880 2.200 18.450 2.600 ;
        RECT  17.720 2.200 17.880 2.610 ;
        RECT  17.360 1.800 17.720 2.610 ;
        RECT  17.260 1.800 17.360 2.600 ;
        RECT  17.050 2.200 17.260 2.600 ;
        END
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.070 1.760 9.470 2.330 ;
        RECT  7.760 1.760 9.070 2.040 ;
        RECT  7.360 1.760 7.760 2.190 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.550 2.110 1.730 2.510 ;
        RECT  1.290 2.110 1.550 3.220 ;
        RECT  0.770 2.920 1.290 3.220 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  18.800 4.640 23.100 5.440 ;
        RECT  18.400 4.480 18.800 5.440 ;
        RECT  17.220 4.640 18.400 5.440 ;
        RECT  16.820 4.480 17.220 5.440 ;
        RECT  15.640 4.640 16.820 5.440 ;
        RECT  14.740 4.480 15.640 5.440 ;
        RECT  10.610 4.640 14.740 5.440 ;
        RECT  10.210 4.480 10.610 5.440 ;
        RECT  9.050 4.640 10.210 5.440 ;
        RECT  8.650 4.480 9.050 5.440 ;
        RECT  1.350 4.640 8.650 5.440 ;
        RECT  0.950 3.980 1.350 5.440 ;
        RECT  0.000 4.640 0.950 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  19.260 -0.400 23.100 0.400 ;
        RECT  18.860 -0.400 19.260 0.560 ;
        RECT  17.680 -0.400 18.860 0.400 ;
        RECT  17.280 -0.400 17.680 0.560 ;
        RECT  16.010 -0.400 17.280 0.400 ;
        RECT  15.850 -0.400 16.010 0.560 ;
        RECT  15.610 -0.400 15.850 1.640 ;
        RECT  10.630 -0.400 15.610 0.400 ;
        RECT  10.230 -0.400 10.630 0.560 ;
        RECT  9.120 -0.400 10.230 0.400 ;
        RECT  8.720 -0.400 9.120 0.560 ;
        RECT  1.350 -0.400 8.720 0.400 ;
        RECT  0.950 -0.400 1.350 0.560 ;
        RECT  0.000 -0.400 0.950 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  22.540 0.640 22.940 1.040 ;
        RECT  22.570 1.440 22.810 4.400 ;
        RECT  22.450 1.440 22.570 1.680 ;
        RECT  20.090 4.160 22.570 4.400 ;
        RECT  21.170 0.640 22.540 0.880 ;
        RECT  22.050 1.280 22.450 1.680 ;
        RECT  21.290 3.000 21.450 3.400 ;
        RECT  21.050 2.460 21.290 3.400 ;
        RECT  20.930 0.640 21.170 2.220 ;
        RECT  20.460 2.460 21.050 2.700 ;
        RECT  19.740 0.640 20.930 0.880 ;
        RECT  20.700 1.820 20.930 2.220 ;
        RECT  20.460 1.130 20.690 1.530 ;
        RECT  20.220 1.130 20.460 2.700 ;
        RECT  18.930 1.280 20.220 1.520 ;
        RECT  19.850 3.420 20.090 4.400 ;
        RECT  18.770 3.420 19.850 3.660 ;
        RECT  19.500 0.640 19.740 1.040 ;
        RECT  19.210 3.900 19.610 4.300 ;
        RECT  16.330 0.800 19.500 1.040 ;
        RECT  6.600 4.000 19.210 4.240 ;
        RECT  18.690 1.280 18.930 3.120 ;
        RECT  18.530 3.420 18.770 3.760 ;
        RECT  18.070 1.280 18.690 1.680 ;
        RECT  18.010 2.880 18.690 3.120 ;
        RECT  8.260 3.520 18.530 3.760 ;
        RECT  17.610 2.880 18.010 3.280 ;
        RECT  16.570 1.280 16.810 2.600 ;
        RECT  16.430 2.360 16.570 2.600 ;
        RECT  16.030 2.360 16.430 3.280 ;
        RECT  16.090 0.800 16.330 2.120 ;
        RECT  15.370 1.880 16.090 2.120 ;
        RECT  14.890 2.360 16.030 2.600 ;
        RECT  15.130 0.640 15.370 2.120 ;
        RECT  13.030 0.640 15.130 0.880 ;
        RECT  14.650 1.120 14.890 2.600 ;
        RECT  13.670 1.120 14.650 1.360 ;
        RECT  13.430 1.120 13.670 3.280 ;
        RECT  13.270 1.120 13.430 1.520 ;
        RECT  10.650 3.040 13.430 3.280 ;
        RECT  13.030 1.760 13.190 2.120 ;
        RECT  12.550 2.400 13.190 2.800 ;
        RECT  12.790 0.640 13.030 2.120 ;
        RECT  12.070 0.700 12.790 0.940 ;
        RECT  12.310 1.180 12.550 2.800 ;
        RECT  11.790 2.560 12.310 2.800 ;
        RECT  11.830 0.700 12.070 2.280 ;
        RECT  11.110 0.700 11.830 0.940 ;
        RECT  11.400 1.870 11.830 2.280 ;
        RECT  11.350 1.180 11.590 1.580 ;
        RECT  11.130 2.560 11.470 2.800 ;
        RECT  11.130 1.340 11.350 1.580 ;
        RECT  10.890 1.340 11.130 2.800 ;
        RECT  10.870 0.700 11.110 1.040 ;
        RECT  6.600 0.800 10.870 1.040 ;
        RECT  10.410 2.020 10.650 3.280 ;
        RECT  10.250 2.020 10.410 2.420 ;
        RECT  9.840 1.280 9.960 2.830 ;
        RECT  9.720 1.280 9.840 3.280 ;
        RECT  9.510 1.280 9.720 1.520 ;
        RECT  9.440 2.590 9.720 3.280 ;
        RECT  8.830 2.590 9.440 2.830 ;
        RECT  8.590 2.280 8.830 2.830 ;
        RECT  8.100 2.280 8.590 2.520 ;
        RECT  7.080 1.280 8.330 1.520 ;
        RECT  7.860 2.860 8.260 3.760 ;
        RECT  7.080 2.860 7.860 3.100 ;
        RECT  6.840 1.280 7.080 3.100 ;
        RECT  6.360 0.800 6.600 1.700 ;
        RECT  5.700 2.020 6.600 2.420 ;
        RECT  6.360 2.740 6.600 4.240 ;
        RECT  5.700 1.300 6.360 1.700 ;
        RECT  5.700 2.740 6.360 3.140 ;
        RECT  4.020 0.660 6.120 0.900 ;
        RECT  5.720 3.510 6.120 4.280 ;
        RECT  4.620 4.040 5.720 4.280 ;
        RECT  4.500 1.460 5.700 1.700 ;
        RECT  4.980 2.180 5.700 2.420 ;
        RECT  5.460 2.900 5.700 3.140 ;
        RECT  5.220 2.900 5.460 3.560 ;
        RECT  4.620 3.320 5.220 3.560 ;
        RECT  4.740 2.180 4.980 2.840 ;
        RECT  4.620 2.600 4.740 2.840 ;
        RECT  2.210 2.600 4.620 3.000 ;
        RECT  3.220 3.320 4.620 3.720 ;
        RECT  3.220 4.040 4.620 4.400 ;
        RECT  4.260 1.460 4.500 2.280 ;
        RECT  3.090 1.880 4.260 2.280 ;
        RECT  3.780 0.660 4.020 1.560 ;
        RECT  3.120 1.160 3.780 1.560 ;
        RECT  2.560 4.120 3.220 4.360 ;
        RECT  2.690 1.240 3.120 1.480 ;
        RECT  2.450 0.800 2.690 1.480 ;
        RECT  2.320 3.470 2.560 4.360 ;
        RECT  0.560 0.800 2.450 1.040 ;
        RECT  0.530 3.470 2.320 3.710 ;
        RECT  1.970 1.280 2.210 3.230 ;
        RECT  1.740 1.280 1.970 1.700 ;
        RECT  1.790 2.830 1.970 3.230 ;
        RECT  1.050 1.460 1.740 1.700 ;
        RECT  0.810 1.460 1.050 2.510 ;
        RECT  0.650 2.110 0.810 2.510 ;
        RECT  0.400 0.770 0.560 1.670 ;
        RECT  0.400 2.820 0.530 4.220 ;
        RECT  0.160 0.770 0.400 4.220 ;
    END
END AFHCINX4

MACRO CMPR32X1
    CLASS CORE ;
    FOREIGN CMPR32X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.850 3.060 13.090 3.460 ;
        RECT  13.090 1.320 13.330 3.460 ;
        RECT  13.330 1.320 13.490 1.720 ;
        RECT  13.330 2.390 13.660 2.650 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.370 2.970 14.720 3.370 ;
        RECT  14.610 1.340 14.720 1.980 ;
        RECT  14.720 1.340 14.980 3.370 ;
        RECT  14.980 1.340 15.010 1.980 ;
        END
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.970 1.960 10.150 2.400 ;
        RECT  10.150 1.960 10.390 4.350 ;
        RECT  10.390 3.950 10.630 4.350 ;
        RECT  10.630 4.060 11.020 4.340 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.210 2.090 ;
        RECT  0.210 1.830 0.460 2.420 ;
        RECT  0.460 2.010 0.570 2.420 ;
        RECT  0.570 2.010 0.810 2.410 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.280 2.320 5.260 2.720 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 4.480 1.390 5.440 ;
        RECT  1.390 4.640 9.470 5.440 ;
        RECT  9.470 4.080 9.870 5.440 ;
        RECT  9.870 4.640 13.610 5.440 ;
        RECT  13.610 3.020 14.010 5.440 ;
        RECT  14.010 4.640 15.180 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        RECT  0.990 -0.400 1.390 0.560 ;
        RECT  1.390 -0.400 4.890 0.400 ;
        RECT  4.890 -0.400 5.290 0.850 ;
        RECT  5.290 -0.400 10.570 0.400 ;
        RECT  10.570 -0.400 10.970 0.560 ;
        RECT  10.970 -0.400 13.850 0.400 ;
        RECT  13.850 -0.400 14.250 1.670 ;
        RECT  14.250 -0.400 15.180 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.930 3.850 13.330 4.250 ;
        RECT  11.750 3.870 12.930 4.110 ;
        RECT  12.510 0.710 12.760 1.110 ;
        RECT  12.270 0.710 12.510 3.590 ;
        RECT  10.330 0.870 12.270 1.110 ;
        RECT  12.110 3.190 12.270 3.590 ;
        RECT  11.750 1.420 11.910 1.820 ;
        RECT  11.510 1.420 11.750 4.110 ;
        RECT  11.350 3.200 11.510 3.600 ;
        RECT  10.710 1.420 10.950 3.510 ;
        RECT  9.850 1.420 10.710 1.660 ;
        RECT  10.670 3.110 10.710 3.510 ;
        RECT  10.090 0.680 10.330 1.110 ;
        RECT  6.610 0.680 10.090 0.920 ;
        RECT  9.610 1.200 9.850 1.660 ;
        RECT  9.370 2.320 9.650 3.610 ;
        RECT  7.200 1.200 9.610 1.440 ;
        RECT  9.250 1.720 9.370 3.610 ;
        RECT  9.130 1.720 9.250 2.640 ;
        RECT  8.370 1.720 8.610 4.360 ;
        RECT  8.090 3.960 8.370 4.360 ;
        RECT  7.850 1.880 8.090 3.430 ;
        RECT  7.730 1.880 7.850 2.120 ;
        RECT  7.450 3.190 7.850 3.430 ;
        RECT  7.490 1.720 7.730 2.120 ;
        RECT  7.430 2.510 7.570 2.910 ;
        RECT  7.290 3.190 7.450 3.590 ;
        RECT  7.200 2.500 7.430 2.910 ;
        RECT  7.050 3.190 7.290 4.360 ;
        RECT  6.960 1.200 7.200 2.910 ;
        RECT  5.820 4.050 7.050 4.360 ;
        RECT  6.690 2.670 6.960 2.910 ;
        RECT  6.530 2.670 6.690 3.510 ;
        RECT  5.870 1.930 6.680 2.330 ;
        RECT  6.370 0.680 6.610 1.590 ;
        RECT  6.450 2.670 6.530 3.770 ;
        RECT  6.290 3.110 6.450 3.770 ;
        RECT  6.210 1.130 6.370 1.590 ;
        RECT  3.770 3.530 6.290 3.770 ;
        RECT  4.610 1.130 6.210 1.370 ;
        RECT  5.870 3.010 5.930 3.250 ;
        RECT  5.630 1.650 5.870 3.250 ;
        RECT  1.910 4.120 5.820 4.360 ;
        RECT  4.090 1.650 5.630 1.890 ;
        RECT  4.050 3.010 5.630 3.250 ;
        RECT  4.370 0.870 4.610 1.370 ;
        RECT  2.690 0.870 4.370 1.110 ;
        RECT  3.850 1.390 4.090 1.890 ;
        RECT  3.530 2.330 3.770 3.770 ;
        RECT  3.470 2.330 3.530 2.570 ;
        RECT  3.230 1.550 3.470 2.570 ;
        RECT  3.010 3.440 3.250 3.840 ;
        RECT  3.210 1.550 3.230 1.790 ;
        RECT  2.970 1.390 3.210 1.790 ;
        RECT  2.950 2.870 3.190 3.110 ;
        RECT  2.430 3.440 3.010 3.680 ;
        RECT  2.710 2.070 2.950 3.110 ;
        RECT  2.690 2.070 2.710 2.310 ;
        RECT  2.450 0.870 2.690 2.310 ;
        RECT  2.190 2.910 2.430 3.680 ;
        RECT  2.170 2.910 2.190 3.310 ;
        RECT  1.930 1.390 2.170 3.310 ;
        RECT  1.840 2.910 1.930 3.310 ;
        RECT  1.670 3.650 1.910 4.360 ;
        RECT  1.470 3.650 1.670 3.890 ;
        RECT  1.470 2.010 1.650 2.410 ;
        RECT  1.230 1.180 1.470 3.890 ;
        RECT  0.570 1.180 1.230 1.420 ;
        RECT  0.170 3.490 1.230 3.890 ;
        RECT  0.170 1.020 0.570 1.420 ;
    END
END CMPR32X1

MACRO CMPR22X1
    CLASS CORE ;
    FOREIGN CMPR22X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 2.950 3.510 3.220 ;
        RECT  3.510 2.950 3.750 3.520 ;
        RECT  3.570 1.190 3.810 1.620 ;
        RECT  3.750 2.950 4.470 3.220 ;
        RECT  3.810 1.380 4.470 1.620 ;
        RECT  4.470 1.380 4.710 3.220 ;
        RECT  4.710 2.950 4.720 3.220 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  7.460 1.270 7.810 1.530 ;
        RECT  7.810 1.260 8.010 1.540 ;
        RECT  8.010 1.230 8.130 1.630 ;
        RECT  8.010 2.970 8.170 3.370 ;
        RECT  8.130 1.230 8.170 1.840 ;
        RECT  8.170 1.230 8.410 3.370 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.840 2.430 2.240 2.830 ;
        RECT  2.240 2.430 2.750 2.750 ;
        RECT  2.750 2.430 2.990 3.220 ;
        RECT  2.990 2.430 3.230 4.250 ;
        RECT  3.230 2.430 3.600 2.670 ;
        RECT  3.600 1.900 3.840 2.670 ;
        RECT  3.840 1.900 4.190 2.140 ;
        RECT  3.230 4.010 5.510 4.250 ;
        RECT  5.510 3.350 5.750 4.250 ;
        RECT  5.750 3.350 6.650 3.590 ;
        RECT  6.650 3.180 6.890 3.590 ;
        RECT  6.890 3.180 7.050 3.580 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.950 1.830 5.850 2.230 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 4.480 1.390 5.440 ;
        RECT  1.390 4.640 6.970 5.440 ;
        RECT  6.970 4.480 7.950 5.440 ;
        RECT  7.950 4.640 8.580 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        RECT  0.990 -0.400 1.390 0.560 ;
        RECT  1.390 -0.400 5.070 0.400 ;
        RECT  5.070 -0.400 5.470 0.560 ;
        RECT  5.470 -0.400 7.900 0.400 ;
        RECT  7.900 -0.400 8.300 0.560 ;
        RECT  8.300 -0.400 8.580 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  7.730 1.950 7.880 2.350 ;
        RECT  7.490 1.950 7.730 4.110 ;
        RECT  7.480 1.950 7.490 2.350 ;
        RECT  6.100 3.870 7.490 4.110 ;
        RECT  7.080 1.960 7.480 2.200 ;
        RECT  6.840 0.640 7.080 2.200 ;
        RECT  6.650 0.640 6.840 0.880 ;
        RECT  6.130 1.310 6.370 3.070 ;
        RECT  5.360 1.310 6.130 1.550 ;
        RECT  5.230 2.830 6.130 3.070 ;
        RECT  5.120 0.860 5.360 1.550 ;
        RECT  4.990 2.830 5.230 3.730 ;
        RECT  4.650 0.860 5.120 1.100 ;
        RECT  4.190 3.490 4.990 3.730 ;
        RECT  4.250 0.670 4.650 1.100 ;
        RECT  3.290 0.670 4.250 0.910 ;
        RECT  3.050 0.670 3.290 2.140 ;
        RECT  1.440 1.900 3.050 2.140 ;
        RECT  2.530 0.700 2.770 1.100 ;
        RECT  2.470 3.640 2.710 4.180 ;
        RECT  0.920 1.380 2.680 1.620 ;
        RECT  0.570 0.860 2.530 1.100 ;
        RECT  0.570 3.940 2.470 4.180 ;
        RECT  1.540 3.380 2.050 3.620 ;
        RECT  1.300 2.980 1.540 3.620 ;
        RECT  1.200 1.900 1.440 2.700 ;
        RECT  0.920 2.980 1.300 3.220 ;
        RECT  0.680 1.380 0.920 3.220 ;
        RECT  0.400 0.700 0.570 1.100 ;
        RECT  0.400 3.500 0.570 4.180 ;
        RECT  0.160 0.700 0.400 4.180 ;
    END
END CMPR22X1

MACRO BENCX2
    CLASS CORE ;
    FOREIGN BENCX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BENCX4 ;
    SIZE 28.380 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN X2
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.360 2.950 17.370 3.210 ;
        RECT  17.370 2.900 17.620 3.210 ;
        RECT  17.620 2.900 19.160 3.140 ;
        RECT  17.370 1.280 19.160 1.520 ;
        RECT  19.160 1.280 19.400 3.140 ;
        RECT  19.400 2.900 19.660 3.140 ;
        END
    END X2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  25.340 0.810 25.420 1.770 ;
        RECT  25.420 0.810 25.740 1.980 ;
        RECT  25.570 2.800 25.970 3.760 ;
        RECT  25.970 2.800 26.780 3.220 ;
        RECT  25.740 1.740 26.780 1.980 ;
        RECT  26.780 0.810 27.010 3.220 ;
        RECT  27.010 0.810 27.180 3.760 ;
        RECT  27.180 2.800 27.410 3.760 ;
        END
    END S
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.510 4.000 12.120 4.240 ;
        RECT  12.120 4.000 12.360 4.400 ;
        RECT  12.360 4.160 13.400 4.400 ;
        RECT  13.400 4.070 13.490 4.400 ;
        RECT  13.490 4.000 13.730 4.400 ;
        RECT  13.730 4.000 21.260 4.240 ;
        END
    END M2
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.440 2.580 6.630 2.820 ;
        RECT  6.630 2.580 6.870 3.760 ;
        RECT  6.870 3.520 8.780 3.760 ;
        RECT  8.780 3.510 8.910 3.770 ;
        RECT  8.910 3.510 9.040 4.250 ;
        RECT  9.040 3.520 9.150 4.250 ;
        RECT  9.150 3.520 9.160 4.170 ;
        RECT  9.160 3.520 12.620 3.760 ;
        RECT  12.620 3.520 12.860 3.920 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.260 2.060 5.390 2.590 ;
        RECT  5.390 2.060 5.830 2.660 ;
        RECT  5.830 2.060 8.020 2.300 ;
        RECT  8.020 0.800 8.260 2.300 ;
        RECT  8.260 0.800 9.420 1.040 ;
        RECT  9.420 0.660 9.660 1.040 ;
        RECT  10.080 2.020 10.500 2.260 ;
        RECT  9.660 0.660 10.500 0.900 ;
        RECT  10.500 0.660 10.740 2.260 ;
        END
    END M0
    PIN A
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.920 0.850 1.320 1.810 ;
        RECT  1.120 2.640 1.430 4.190 ;
        RECT  1.320 1.570 1.430 1.810 ;
        RECT  1.430 2.370 1.520 4.190 ;
        RECT  1.520 2.370 1.530 3.220 ;
        RECT  1.530 2.370 1.640 2.970 ;
        RECT  1.430 1.570 1.640 1.840 ;
        RECT  1.640 1.570 1.880 2.970 ;
        RECT  1.880 1.570 2.370 1.810 ;
        RECT  1.880 2.730 2.430 2.970 ;
        RECT  2.430 2.730 2.650 3.220 ;
        RECT  2.370 0.850 2.770 1.810 ;
        RECT  2.650 2.730 2.890 4.190 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.400 5.440 ;
        RECT  0.400 3.530 0.800 5.440 ;
        RECT  0.800 4.640 1.850 5.440 ;
        RECT  1.850 3.530 2.250 5.440 ;
        RECT  2.250 4.640 3.290 5.440 ;
        RECT  3.290 4.090 3.690 5.440 ;
        RECT  3.690 4.640 4.750 5.440 ;
        RECT  4.750 4.090 5.150 5.440 ;
        RECT  5.150 4.640 6.580 5.440 ;
        RECT  6.580 4.480 6.980 5.440 ;
        RECT  6.980 4.640 8.270 5.440 ;
        RECT  8.270 4.060 8.670 5.440 ;
        RECT  8.670 4.640 10.100 5.440 ;
        RECT  10.100 4.480 10.500 5.440 ;
        RECT  10.500 4.640 11.480 5.440 ;
        RECT  11.480 4.480 11.880 5.440 ;
        RECT  11.880 4.640 15.460 5.440 ;
        RECT  15.460 4.480 15.860 5.440 ;
        RECT  15.860 4.640 16.840 5.440 ;
        RECT  16.840 4.480 17.240 5.440 ;
        RECT  17.240 4.640 18.470 5.440 ;
        RECT  18.470 4.480 18.870 5.440 ;
        RECT  18.870 4.640 20.080 5.440 ;
        RECT  20.080 4.480 20.480 5.440 ;
        RECT  20.480 4.640 21.430 5.440 ;
        RECT  21.430 4.480 21.830 5.440 ;
        RECT  21.830 4.640 23.420 5.440 ;
        RECT  23.420 4.480 23.820 5.440 ;
        RECT  23.820 4.640 24.740 5.440 ;
        RECT  24.740 4.480 24.850 5.440 ;
        RECT  24.850 3.310 25.250 5.440 ;
        RECT  25.250 4.640 26.290 5.440 ;
        RECT  26.290 3.490 26.690 5.440 ;
        RECT  26.690 4.640 27.730 5.440 ;
        RECT  27.730 2.740 28.130 5.440 ;
        RECT  28.130 4.640 28.380 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.190 0.400 ;
        RECT  0.190 -0.400 0.590 1.620 ;
        RECT  0.590 -0.400 1.640 0.400 ;
        RECT  1.640 -0.400 2.040 1.060 ;
        RECT  2.040 -0.400 3.170 0.400 ;
        RECT  3.170 -0.400 3.570 0.560 ;
        RECT  3.570 -0.400 4.580 0.400 ;
        RECT  4.580 -0.400 4.980 0.560 ;
        RECT  4.980 -0.400 6.220 0.400 ;
        RECT  6.220 -0.400 6.620 0.560 ;
        RECT  6.620 -0.400 8.690 0.400 ;
        RECT  8.690 -0.400 9.090 0.560 ;
        RECT  9.090 -0.400 11.780 0.400 ;
        RECT  11.780 -0.400 12.180 0.560 ;
        RECT  12.180 -0.400 15.510 0.400 ;
        RECT  15.510 -0.400 15.910 0.560 ;
        RECT  15.910 -0.400 16.580 0.400 ;
        RECT  16.580 -0.400 16.980 0.560 ;
        RECT  16.980 -0.400 18.180 0.400 ;
        RECT  18.180 -0.400 18.580 0.560 ;
        RECT  18.580 -0.400 19.780 0.400 ;
        RECT  19.780 -0.400 20.180 0.560 ;
        RECT  20.180 -0.400 21.560 0.400 ;
        RECT  21.560 -0.400 21.960 0.560 ;
        RECT  21.960 -0.400 23.170 0.400 ;
        RECT  23.170 -0.400 23.570 0.560 ;
        RECT  23.570 -0.400 24.540 0.400 ;
        RECT  24.540 -0.400 24.940 0.560 ;
        RECT  24.940 -0.400 26.140 0.400 ;
        RECT  26.140 -0.400 26.380 1.300 ;
        RECT  26.380 -0.400 27.580 0.400 ;
        RECT  27.580 -0.400 27.820 1.770 ;
        RECT  27.820 -0.400 28.380 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  25.230 2.270 26.520 2.510 ;
        RECT  24.990 2.270 25.230 3.070 ;
        RECT  24.970 2.270 24.990 2.510 ;
        RECT  24.310 2.830 24.990 3.070 ;
        RECT  24.730 1.450 24.970 2.510 ;
        RECT  23.870 1.450 24.730 1.690 ;
        RECT  24.070 2.830 24.310 3.790 ;
        RECT  23.710 2.090 24.110 2.490 ;
        RECT  23.460 2.100 23.710 2.490 ;
        RECT  23.220 1.660 23.460 3.660 ;
        RECT  21.820 1.660 23.220 1.900 ;
        RECT  20.630 3.420 23.220 3.660 ;
        RECT  22.390 1.080 22.770 1.320 ;
        RECT  22.530 2.160 22.770 2.970 ;
        RECT  19.890 2.160 22.530 2.400 ;
        RECT  22.150 0.880 22.390 1.320 ;
        RECT  20.780 0.880 22.150 1.120 ;
        RECT  20.190 2.660 22.130 2.900 ;
        RECT  21.580 1.390 21.820 1.900 ;
        RECT  21.040 1.390 21.580 1.630 ;
        RECT  20.540 0.880 20.780 1.420 ;
        RECT  20.320 1.180 20.540 1.420 ;
        RECT  19.950 2.660 20.190 3.760 ;
        RECT  15.630 3.520 19.950 3.760 ;
        RECT  19.650 0.800 19.890 2.400 ;
        RECT  15.140 0.800 19.650 1.040 ;
        RECT  16.770 2.090 18.900 2.330 ;
        RECT  16.550 1.380 16.770 2.330 ;
        RECT  16.530 1.380 16.550 3.230 ;
        RECT  15.790 1.380 16.530 1.620 ;
        RECT  16.310 2.090 16.530 3.230 ;
        RECT  15.390 2.280 15.630 3.760 ;
        RECT  15.070 0.640 15.140 1.040 ;
        RECT  15.020 0.640 15.070 2.510 ;
        RECT  14.830 0.640 15.020 3.490 ;
        RECT  12.740 0.640 14.830 0.880 ;
        RECT  14.780 2.270 14.830 3.490 ;
        RECT  14.540 1.120 14.590 2.020 ;
        RECT  14.350 1.120 14.540 3.710 ;
        RECT  13.360 1.120 14.350 1.360 ;
        RECT  14.300 1.700 14.350 3.710 ;
        RECT  13.840 3.470 14.300 3.710 ;
        RECT  13.820 1.710 14.060 3.230 ;
        RECT  13.040 1.710 13.820 1.950 ;
        RECT  12.210 2.990 13.820 3.230 ;
        RECT  13.340 2.220 13.580 2.630 ;
        RECT  11.940 2.390 13.340 2.630 ;
        RECT  12.800 1.280 13.040 1.950 ;
        RECT  12.640 1.280 12.800 1.520 ;
        RECT  12.500 0.640 12.740 1.040 ;
        RECT  12.380 1.870 12.540 2.110 ;
        RECT  12.380 0.800 12.500 1.040 ;
        RECT  12.140 0.800 12.380 2.110 ;
        RECT  11.510 1.870 12.140 2.110 ;
        RECT  11.700 2.390 11.940 3.280 ;
        RECT  9.510 3.040 11.700 3.280 ;
        RECT  11.310 1.180 11.510 2.110 ;
        RECT  11.270 1.180 11.310 2.800 ;
        RECT  11.070 1.870 11.270 2.800 ;
        RECT  10.690 2.560 11.070 2.800 ;
        RECT  9.950 1.180 10.190 1.680 ;
        RECT  9.500 1.440 9.950 1.680 ;
        RECT  9.500 2.910 9.510 3.280 ;
        RECT  9.270 1.440 9.500 3.280 ;
        RECT  9.260 1.440 9.270 3.150 ;
        RECT  9.070 2.910 9.260 3.150 ;
        RECT  8.500 1.280 8.740 3.260 ;
        RECT  7.140 3.020 8.500 3.260 ;
        RECT  7.540 1.230 7.780 1.790 ;
        RECT  6.230 4.000 7.770 4.240 ;
        RECT  4.920 1.550 7.540 1.790 ;
        RECT  5.410 1.050 7.140 1.290 ;
        RECT  5.990 3.120 6.230 4.240 ;
        RECT  4.920 3.120 5.990 3.360 ;
        RECT  4.680 1.550 4.920 3.360 ;
        RECT  3.700 2.070 4.680 2.470 ;
        RECT  3.370 3.610 4.420 3.850 ;
        RECT  3.370 1.140 4.250 1.380 ;
        RECT  3.130 1.140 3.370 3.850 ;
        RECT  2.130 2.150 3.130 2.390 ;
    END
END BENCX2

MACRO BENCX1
    CLASS CORE ;
    FOREIGN BENCX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BENCX4 ;
    SIZE 21.120 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN X2
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.060 2.950 14.190 3.210 ;
        RECT  14.190 2.900 14.320 3.210 ;
        RECT  14.320 2.900 14.380 3.200 ;
        RECT  13.710 1.280 14.380 1.520 ;
        RECT  14.380 1.280 14.500 3.200 ;
        RECT  14.500 1.280 14.620 3.140 ;
        END
    END X2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  19.750 2.800 20.110 3.760 ;
        RECT  19.820 0.810 20.110 1.770 ;
        RECT  20.110 0.810 20.150 3.760 ;
        RECT  20.150 0.810 20.220 3.270 ;
        RECT  20.220 1.320 20.350 3.270 ;
        RECT  20.350 2.950 20.370 3.270 ;
        END
    END S
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.970 4.000 7.460 4.240 ;
        RECT  7.460 4.000 7.720 4.330 ;
        RECT  7.720 4.000 8.870 4.240 ;
        RECT  8.870 4.000 9.110 4.400 ;
        RECT  9.110 4.160 11.010 4.400 ;
        RECT  11.010 4.000 11.430 4.400 ;
        RECT  11.430 4.000 16.120 4.240 ;
        END
    END M2
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.900 2.750 4.090 2.990 ;
        RECT  4.090 2.750 4.330 3.760 ;
        RECT  4.330 3.520 6.140 3.760 ;
        RECT  6.140 3.510 6.290 3.770 ;
        RECT  6.290 3.510 6.400 3.820 ;
        RECT  6.400 3.520 6.690 3.820 ;
        RECT  6.690 3.520 9.350 3.760 ;
        RECT  9.350 3.520 9.590 3.920 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.390 2.980 2.650 ;
        RECT  2.980 2.270 3.100 2.650 ;
        RECT  3.100 2.270 3.220 2.640 ;
        RECT  3.220 2.270 5.480 2.510 ;
        RECT  5.480 0.800 5.720 2.510 ;
        RECT  5.720 0.800 6.890 1.040 ;
        RECT  6.890 0.640 7.130 1.040 ;
        RECT  7.130 0.640 7.920 0.880 ;
        END
    END M0
    PIN A
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.320 1.590 0.560 2.970 ;
        RECT  0.560 1.590 0.770 1.830 ;
        RECT  0.560 2.730 0.860 2.970 ;
        RECT  0.860 2.730 0.990 3.210 ;
        RECT  0.770 1.410 1.120 1.830 ;
        RECT  1.120 1.410 1.200 1.810 ;
        RECT  0.990 2.730 1.230 4.190 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.190 5.440 ;
        RECT  0.190 3.530 0.590 5.440 ;
        RECT  0.590 4.640 1.630 5.440 ;
        RECT  1.630 4.090 2.030 5.440 ;
        RECT  2.030 4.640 4.040 5.440 ;
        RECT  4.040 4.480 4.440 5.440 ;
        RECT  4.440 4.640 5.740 5.440 ;
        RECT  5.740 4.060 6.140 5.440 ;
        RECT  6.140 4.640 8.210 5.440 ;
        RECT  8.210 4.480 8.610 5.440 ;
        RECT  8.610 4.640 13.400 5.440 ;
        RECT  13.400 4.480 13.800 5.440 ;
        RECT  13.800 4.640 14.980 5.440 ;
        RECT  14.980 4.480 15.380 5.440 ;
        RECT  15.380 4.640 16.280 5.440 ;
        RECT  16.280 4.480 16.680 5.440 ;
        RECT  16.680 4.640 18.950 5.440 ;
        RECT  18.950 4.480 19.030 5.440 ;
        RECT  19.030 3.310 19.430 5.440 ;
        RECT  19.430 4.640 20.550 5.440 ;
        RECT  20.550 3.490 20.790 5.440 ;
        RECT  20.790 4.640 21.120 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 1.080 ;
        RECT  0.560 -0.400 1.510 0.400 ;
        RECT  1.510 -0.400 1.910 0.560 ;
        RECT  1.910 -0.400 2.710 0.400 ;
        RECT  2.710 -0.400 3.110 0.560 ;
        RECT  3.110 -0.400 6.150 0.400 ;
        RECT  6.150 -0.400 6.550 0.560 ;
        RECT  6.550 -0.400 8.890 0.400 ;
        RECT  8.890 -0.400 9.290 0.560 ;
        RECT  9.290 -0.400 12.920 0.400 ;
        RECT  12.920 -0.400 13.320 0.560 ;
        RECT  13.320 -0.400 14.520 0.400 ;
        RECT  14.520 -0.400 14.920 0.560 ;
        RECT  14.920 -0.400 16.540 0.400 ;
        RECT  16.540 -0.400 16.940 0.560 ;
        RECT  16.940 -0.400 17.730 0.400 ;
        RECT  17.730 -0.400 18.130 0.560 ;
        RECT  18.130 -0.400 19.020 0.400 ;
        RECT  19.020 -0.400 19.420 0.560 ;
        RECT  19.420 -0.400 20.620 0.400 ;
        RECT  20.620 -0.400 20.860 1.740 ;
        RECT  20.860 -0.400 21.120 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  19.410 2.070 19.860 2.470 ;
        RECT  19.170 1.450 19.410 3.070 ;
        RECT  18.350 1.450 19.170 1.690 ;
        RECT  18.490 2.830 19.170 3.070 ;
        RECT  17.910 2.090 18.730 2.490 ;
        RECT  18.250 2.830 18.490 3.790 ;
        RECT  17.710 2.090 17.910 3.660 ;
        RECT  17.670 1.560 17.710 3.660 ;
        RECT  17.470 1.560 17.670 2.330 ;
        RECT  15.420 3.420 17.670 3.660 ;
        RECT  15.820 1.560 17.470 1.800 ;
        RECT  16.300 1.080 17.440 1.320 ;
        RECT  15.130 2.120 17.230 2.360 ;
        RECT  15.140 2.800 16.900 3.040 ;
        RECT  16.060 0.640 16.300 1.320 ;
        RECT  15.420 0.640 16.060 0.880 ;
        RECT  15.580 1.360 15.820 1.800 ;
        RECT  15.420 1.360 15.580 1.600 ;
        RECT  14.900 2.800 15.140 3.760 ;
        RECT  14.890 0.800 15.130 2.360 ;
        RECT  12.450 3.520 14.900 3.760 ;
        RECT  12.040 0.800 14.890 1.040 ;
        RECT  12.930 2.090 13.930 2.330 ;
        RECT  12.690 1.450 12.930 3.280 ;
        RECT  12.450 1.450 12.690 1.690 ;
        RECT  12.210 1.280 12.450 1.690 ;
        RECT  12.210 2.300 12.450 3.760 ;
        RECT  11.970 0.640 12.040 1.040 ;
        RECT  11.730 0.640 11.970 3.610 ;
        RECT  9.870 0.640 11.730 0.880 ;
        RECT  11.250 1.120 11.490 3.520 ;
        RECT  10.260 1.120 11.250 1.360 ;
        RECT  10.570 3.280 11.250 3.520 ;
        RECT  10.770 1.830 11.010 3.030 ;
        RECT  10.010 1.830 10.770 2.070 ;
        RECT  10.270 2.790 10.770 3.030 ;
        RECT  8.400 2.310 10.530 2.550 ;
        RECT  10.030 2.790 10.270 3.270 ;
        RECT  8.940 3.030 10.030 3.270 ;
        RECT  9.770 1.280 10.010 2.070 ;
        RECT  9.630 0.640 9.870 1.040 ;
        RECT  9.480 1.280 9.770 1.520 ;
        RECT  9.070 0.800 9.630 1.040 ;
        RECT  9.070 1.830 9.430 2.070 ;
        RECT  8.830 0.800 9.070 2.070 ;
        RECT  8.760 1.260 8.830 2.070 ;
        RECT  8.120 1.260 8.760 1.500 ;
        RECT  7.920 1.830 8.760 2.070 ;
        RECT  8.160 2.310 8.400 3.280 ;
        RECT  6.970 3.040 8.160 3.280 ;
        RECT  7.680 1.830 7.920 2.800 ;
        RECT  7.620 1.260 7.800 1.500 ;
        RECT  7.410 2.560 7.680 2.800 ;
        RECT  7.380 1.260 7.620 1.580 ;
        RECT  6.960 1.340 7.380 1.580 ;
        RECT  6.960 3.020 6.970 3.280 ;
        RECT  6.730 1.340 6.960 3.280 ;
        RECT  6.720 1.340 6.730 3.260 ;
        RECT  6.530 3.020 6.720 3.260 ;
        RECT  5.960 1.280 6.200 3.260 ;
        RECT  4.600 3.020 5.960 3.260 ;
        RECT  3.690 4.000 5.300 4.240 ;
        RECT  5.000 0.910 5.240 1.340 ;
        RECT  5.000 1.620 5.240 2.030 ;
        RECT  3.500 1.100 5.000 1.340 ;
        RECT  2.190 1.620 5.000 1.860 ;
        RECT  3.450 3.430 3.690 4.240 ;
        RECT  3.030 3.430 3.450 3.670 ;
        RECT  2.790 3.060 3.030 3.670 ;
        RECT  2.190 3.060 2.790 3.300 ;
        RECT  2.530 4.150 2.760 4.390 ;
        RECT  1.710 1.140 2.590 1.380 ;
        RECT  2.290 3.610 2.530 4.390 ;
        RECT  1.710 3.610 2.290 3.850 ;
        RECT  1.950 1.620 2.190 3.300 ;
        RECT  1.470 1.140 1.710 3.850 ;
        RECT  0.800 2.150 1.470 2.390 ;
    END
END BENCX1

MACRO XOR2XL
    CLASS CORE ;
    FOREIGN XOR2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 2.940 4.830 3.540 ;
        RECT  4.720 1.100 4.830 1.500 ;
        RECT  4.830 1.100 5.070 3.540 ;
        RECT  5.070 1.100 5.120 1.500 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 1.000 3.210 ;
        RECT  1.000 2.410 1.120 3.210 ;
        RECT  1.120 2.410 1.240 3.200 ;
        RECT  1.240 2.410 1.400 2.650 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.610 1.650 0.850 2.090 ;
        RECT  0.850 1.840 0.870 2.090 ;
        RECT  0.870 1.850 1.520 2.090 ;
        RECT  1.520 1.830 1.780 2.090 ;
        RECT  1.780 1.850 1.870 2.090 ;
        RECT  1.870 1.850 2.110 2.480 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.560 5.440 ;
        RECT  0.560 4.480 0.960 5.440 ;
        RECT  0.960 4.640 4.080 5.440 ;
        RECT  4.080 4.480 4.480 5.440 ;
        RECT  4.480 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.550 0.400 ;
        RECT  0.550 -0.400 0.950 0.560 ;
        RECT  0.950 -0.400 4.060 0.400 ;
        RECT  4.060 -0.400 4.460 0.560 ;
        RECT  4.460 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.330 1.740 4.570 2.140 ;
        RECT  4.170 1.740 4.330 1.980 ;
        RECT  3.930 0.800 4.170 1.980 ;
        RECT  3.070 0.800 3.930 1.040 ;
        RECT  3.560 3.530 3.800 3.930 ;
        RECT  3.550 1.280 3.590 1.680 ;
        RECT  2.000 3.680 3.560 3.920 ;
        RECT  3.310 1.280 3.550 3.290 ;
        RECT  2.830 0.800 3.070 3.440 ;
        RECT  1.440 4.160 3.040 4.400 ;
        RECT  2.800 0.800 2.830 1.100 ;
        RECT  2.410 3.200 2.830 3.440 ;
        RECT  2.560 0.700 2.800 1.100 ;
        RECT  2.350 1.340 2.590 2.960 ;
        RECT  2.090 1.340 2.350 1.580 ;
        RECT  2.000 2.720 2.350 2.960 ;
        RECT  1.430 0.640 2.240 0.880 ;
        RECT  1.850 1.220 2.090 1.580 ;
        RECT  1.760 2.720 2.000 3.920 ;
        RECT  1.690 1.220 1.850 1.460 ;
        RECT  1.200 3.680 1.440 4.400 ;
        RECT  1.190 0.640 1.430 1.100 ;
        RECT  0.480 3.680 1.200 3.920 ;
        RECT  0.560 0.860 1.190 1.100 ;
        RECT  0.370 0.860 0.560 1.320 ;
        RECT  0.370 3.520 0.480 3.920 ;
        RECT  0.320 0.860 0.370 3.920 ;
        RECT  0.240 1.080 0.320 3.920 ;
        RECT  0.130 1.080 0.240 3.790 ;
    END
END XOR2XL

MACRO XOR2X4
    CLASS CORE ;
    FOREIGN XOR2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ XOR2XL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  10.670 2.940 10.680 4.340 ;
        RECT  10.480 1.380 10.680 1.780 ;
        RECT  10.680 2.890 10.920 4.340 ;
        RECT  10.680 1.370 10.920 1.790 ;
        RECT  10.920 1.370 11.110 4.340 ;
        RECT  11.110 1.370 11.340 3.640 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.540 2.070 1.520 2.470 ;
        RECT  1.520 2.070 1.780 2.650 ;
        RECT  1.780 2.070 2.040 2.470 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.130 2.170 7.460 2.570 ;
        RECT  7.460 2.170 7.530 2.650 ;
        RECT  7.530 2.250 7.710 2.650 ;
        RECT  7.710 2.390 7.720 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.180 5.440 ;
        RECT  0.180 4.010 0.580 5.440 ;
        RECT  0.580 4.640 1.570 5.440 ;
        RECT  1.570 4.130 1.970 5.440 ;
        RECT  1.970 4.640 3.050 5.440 ;
        RECT  3.050 4.210 3.450 5.440 ;
        RECT  3.450 4.640 8.390 5.440 ;
        RECT  8.390 4.480 8.790 5.440 ;
        RECT  8.790 4.640 9.880 5.440 ;
        RECT  9.880 4.150 10.120 5.440 ;
        RECT  10.120 4.640 11.390 5.440 ;
        RECT  11.390 4.150 11.630 5.440 ;
        RECT  11.630 4.640 11.880 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.420 0.400 ;
        RECT  0.420 -0.400 0.430 0.850 ;
        RECT  0.430 -0.400 0.830 1.050 ;
        RECT  0.830 -0.400 0.840 0.850 ;
        RECT  0.840 -0.400 1.760 0.400 ;
        RECT  1.760 -0.400 1.770 0.850 ;
        RECT  1.770 -0.400 2.170 1.050 ;
        RECT  2.170 -0.400 2.180 0.850 ;
        RECT  2.180 -0.400 3.110 0.400 ;
        RECT  3.110 -0.400 3.510 0.560 ;
        RECT  3.510 -0.400 8.370 0.400 ;
        RECT  8.370 -0.400 8.770 0.560 ;
        RECT  8.770 -0.400 9.750 0.400 ;
        RECT  9.750 -0.400 10.150 0.560 ;
        RECT  10.150 -0.400 11.080 0.400 ;
        RECT  11.080 -0.400 11.090 0.780 ;
        RECT  11.090 -0.400 11.490 0.980 ;
        RECT  11.490 -0.400 11.500 0.780 ;
        RECT  11.500 -0.400 11.880 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.240 2.180 10.640 2.580 ;
        RECT  10.200 2.180 10.240 2.420 ;
        RECT  9.960 0.860 10.200 2.420 ;
        RECT  8.040 0.860 9.960 1.100 ;
        RECT  9.290 1.380 9.530 3.410 ;
        RECT  9.080 1.380 9.290 1.890 ;
        RECT  9.070 3.010 9.290 3.410 ;
        RECT  7.280 1.650 9.080 1.890 ;
        RECT  8.760 2.300 8.970 2.700 ;
        RECT  8.520 2.300 8.760 4.170 ;
        RECT  7.290 3.930 8.520 4.170 ;
        RECT  7.960 0.860 8.040 1.280 ;
        RECT  7.630 3.250 8.030 3.650 ;
        RECT  7.640 0.790 7.960 1.280 ;
        RECT  6.520 0.790 7.640 1.030 ;
        RECT  6.530 3.250 7.630 3.490 ;
        RECT  7.210 3.770 7.290 4.170 ;
        RECT  6.880 1.310 7.280 1.890 ;
        RECT  6.890 3.770 7.210 4.250 ;
        RECT  3.990 4.010 6.890 4.250 ;
        RECT  6.850 1.650 6.880 1.890 ;
        RECT  6.610 1.650 6.850 2.970 ;
        RECT  5.770 2.730 6.610 2.970 ;
        RECT  6.130 3.250 6.530 3.730 ;
        RECT  6.330 0.790 6.520 1.360 ;
        RECT  6.090 0.790 6.330 1.830 ;
        RECT  5.090 3.490 6.130 3.730 ;
        RECT  5.090 1.590 6.090 1.830 ;
        RECT  5.370 2.730 5.770 3.210 ;
        RECT  5.360 0.860 5.760 1.310 ;
        RECT  2.840 0.860 5.360 1.100 ;
        RECT  5.000 1.590 5.090 3.730 ;
        RECT  4.850 1.450 5.000 3.730 ;
        RECT  4.600 1.450 4.850 1.830 ;
        RECT  4.610 3.320 4.850 3.730 ;
        RECT  4.270 2.150 4.570 2.560 ;
        RECT  4.030 1.390 4.270 3.390 ;
        RECT  3.860 1.390 4.030 1.790 ;
        RECT  3.870 2.990 4.030 3.390 ;
        RECT  3.750 3.680 3.990 4.250 ;
        RECT  2.790 3.680 3.750 3.920 ;
        RECT  2.790 0.860 2.840 3.330 ;
        RECT  2.600 0.860 2.790 3.920 ;
        RECT  2.440 1.390 2.600 1.790 ;
        RECT  2.550 3.010 2.600 3.920 ;
        RECT  0.850 3.010 2.550 3.410 ;
        RECT  1.500 1.470 2.440 1.710 ;
        RECT  1.100 1.390 1.500 1.790 ;
    END
END XOR2X4

MACRO XOR2X2
    CLASS CORE ;
    FOREIGN XOR2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ XOR2XL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.050 2.940 6.220 4.340 ;
        RECT  6.220 2.740 6.490 4.340 ;
        RECT  6.490 2.740 6.550 4.140 ;
        RECT  6.270 0.800 6.550 1.540 ;
        RECT  6.550 0.800 6.620 4.140 ;
        RECT  6.620 0.800 6.670 3.190 ;
        RECT  6.670 1.300 6.790 3.190 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 0.980 3.210 ;
        RECT  0.980 2.680 1.220 3.210 ;
        RECT  1.220 2.680 1.320 2.920 ;
        RECT  1.320 2.420 1.560 2.920 ;
        RECT  1.560 2.420 1.850 2.660 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 1.900 0.920 2.300 ;
        RECT  0.920 1.900 2.100 2.140 ;
        RECT  2.100 1.900 2.340 2.650 ;
        RECT  2.340 2.220 2.520 2.650 ;
        RECT  2.520 2.220 3.280 2.460 ;
        RECT  3.280 2.060 3.520 2.460 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.820 5.440 ;
        RECT  0.820 3.660 1.060 5.440 ;
        RECT  1.060 4.640 2.270 5.440 ;
        RECT  2.270 3.730 2.670 5.440 ;
        RECT  2.670 4.640 5.560 5.440 ;
        RECT  5.560 3.870 5.800 5.440 ;
        RECT  5.800 4.640 7.260 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 2.440 0.400 ;
        RECT  2.440 -0.400 2.840 0.560 ;
        RECT  2.840 -0.400 5.440 0.400 ;
        RECT  5.440 -0.400 5.840 0.560 ;
        RECT  5.840 -0.400 7.260 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.070 1.780 6.310 2.350 ;
        RECT  5.580 1.780 6.070 2.020 ;
        RECT  5.460 2.260 5.620 2.500 ;
        RECT  5.340 0.870 5.580 2.020 ;
        RECT  5.220 2.260 5.460 3.620 ;
        RECT  4.480 0.870 5.340 1.110 ;
        RECT  4.960 3.380 5.220 3.620 ;
        RECT  4.720 1.380 4.960 3.140 ;
        RECT  4.720 3.380 4.960 4.180 ;
        RECT  3.430 3.940 4.720 4.180 ;
        RECT  4.240 0.870 4.480 3.500 ;
        RECT  3.880 0.870 4.240 1.270 ;
        RECT  4.150 3.260 4.240 3.500 ;
        RECT  3.750 3.260 4.150 3.660 ;
        RECT  3.760 1.540 4.000 2.980 ;
        RECT  3.620 1.540 3.760 1.780 ;
        RECT  3.430 2.740 3.760 2.980 ;
        RECT  3.380 0.690 3.620 1.780 ;
        RECT  3.190 2.740 3.430 4.180 ;
        RECT  3.160 0.690 3.380 1.100 ;
        RECT  3.110 2.990 3.190 4.180 ;
        RECT  1.630 0.860 3.160 1.100 ;
        RECT  0.570 1.380 3.140 1.620 ;
        RECT  3.030 2.990 3.110 3.970 ;
        RECT  1.910 3.210 3.030 3.450 ;
        RECT  1.510 3.210 1.910 4.110 ;
        RECT  0.400 1.230 0.570 1.620 ;
        RECT  0.490 3.000 0.520 4.400 ;
        RECT  0.400 2.840 0.490 4.400 ;
        RECT  0.280 1.230 0.400 4.400 ;
        RECT  0.250 1.230 0.280 3.240 ;
        RECT  0.160 1.230 0.250 3.080 ;
    END
END XOR2X2

MACRO XOR2X1
    CLASS CORE ;
    FOREIGN XOR2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ XOR2XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 2.940 4.830 3.540 ;
        RECT  4.670 1.100 4.830 1.500 ;
        RECT  4.830 1.100 5.070 3.540 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 1.000 3.210 ;
        RECT  1.000 2.410 1.120 3.210 ;
        RECT  1.120 2.410 1.240 3.200 ;
        RECT  1.240 2.410 1.400 2.650 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.610 1.600 0.850 2.090 ;
        RECT  0.850 1.840 0.870 2.090 ;
        RECT  0.870 1.850 1.520 2.090 ;
        RECT  1.520 1.830 1.780 2.090 ;
        RECT  1.780 1.850 1.860 2.090 ;
        RECT  1.860 1.850 2.100 2.480 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.560 5.440 ;
        RECT  0.560 4.480 0.960 5.440 ;
        RECT  0.960 4.640 4.080 5.440 ;
        RECT  4.080 4.480 4.480 5.440 ;
        RECT  4.480 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.660 0.400 ;
        RECT  0.660 -0.400 1.060 0.560 ;
        RECT  1.060 -0.400 4.330 0.400 ;
        RECT  4.330 -0.400 4.730 0.560 ;
        RECT  4.730 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.320 1.740 4.560 2.140 ;
        RECT  4.090 1.740 4.320 1.980 ;
        RECT  3.850 0.720 4.090 1.980 ;
        RECT  3.060 0.720 3.850 0.960 ;
        RECT  3.670 3.700 3.830 4.100 ;
        RECT  3.430 3.680 3.670 4.100 ;
        RECT  3.540 1.200 3.610 1.600 ;
        RECT  3.370 1.200 3.540 3.280 ;
        RECT  1.920 3.680 3.430 3.920 ;
        RECT  3.300 1.360 3.370 3.280 ;
        RECT  2.820 0.720 3.060 3.440 ;
        RECT  1.440 4.160 3.040 4.400 ;
        RECT  2.580 0.700 2.820 1.100 ;
        RECT  2.390 3.200 2.820 3.440 ;
        RECT  2.340 1.340 2.580 2.960 ;
        RECT  1.540 0.640 2.340 0.880 ;
        RECT  1.590 1.340 2.340 1.580 ;
        RECT  1.920 2.720 2.340 2.960 ;
        RECT  1.680 2.720 1.920 3.920 ;
        RECT  1.300 0.640 1.540 1.100 ;
        RECT  1.200 3.680 1.440 4.400 ;
        RECT  0.570 0.860 1.300 1.100 ;
        RECT  0.490 3.680 1.200 3.920 ;
        RECT  0.370 0.860 0.570 1.320 ;
        RECT  0.370 3.520 0.490 3.920 ;
        RECT  0.330 0.860 0.370 3.920 ;
        RECT  0.250 1.080 0.330 3.920 ;
        RECT  0.130 1.080 0.250 3.790 ;
    END
END XOR2X1

MACRO XNOR2XL
    CLASS CORE ;
    FOREIGN XNOR2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.820 2.950 4.950 3.210 ;
        RECT  4.950 2.950 5.100 3.260 ;
        RECT  5.100 2.860 5.370 3.260 ;
        RECT  5.370 1.400 5.500 3.260 ;
        RECT  5.500 1.400 5.610 3.100 ;
        RECT  5.610 1.400 5.770 1.840 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.470 2.180 1.870 2.660 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.760 2.100 0.770 2.500 ;
        RECT  0.770 1.820 1.120 2.510 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.670 5.440 ;
        RECT  0.670 3.860 0.680 5.440 ;
        RECT  0.680 3.660 1.080 5.440 ;
        RECT  1.080 3.860 1.090 5.440 ;
        RECT  1.090 4.640 4.280 5.440 ;
        RECT  4.280 4.480 4.680 5.440 ;
        RECT  4.680 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.530 0.400 ;
        RECT  0.530 -0.400 0.930 0.560 ;
        RECT  0.930 -0.400 4.360 0.400 ;
        RECT  4.360 -0.400 4.760 0.560 ;
        RECT  4.760 -0.400 5.940 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.930 1.960 5.130 2.360 ;
        RECT  4.730 0.860 4.930 2.360 ;
        RECT  4.690 0.860 4.730 2.200 ;
        RECT  3.080 0.860 4.690 1.100 ;
        RECT  3.640 3.510 4.040 4.120 ;
        RECT  3.740 1.380 3.840 1.780 ;
        RECT  3.500 1.380 3.740 3.230 ;
        RECT  2.380 3.510 3.640 3.750 ;
        RECT  3.440 1.380 3.500 1.780 ;
        RECT  3.340 2.830 3.500 3.230 ;
        RECT  3.000 0.860 3.080 1.770 ;
        RECT  2.840 0.860 3.000 3.230 ;
        RECT  2.760 1.370 2.840 3.230 ;
        RECT  2.680 1.370 2.760 1.770 ;
        RECT  2.660 2.830 2.760 3.230 ;
        RECT  1.600 4.030 2.720 4.270 ;
        RECT  2.140 1.390 2.380 3.750 ;
        RECT  2.000 1.390 2.140 1.790 ;
        RECT  1.880 3.020 2.140 3.420 ;
        RECT  1.760 0.670 2.120 0.910 ;
        RECT  1.520 0.670 1.760 1.550 ;
        RECT  1.360 3.140 1.600 4.270 ;
        RECT  0.490 1.310 1.520 1.550 ;
        RECT  0.570 3.140 1.360 3.380 ;
        RECT  0.410 2.770 0.570 3.380 ;
        RECT  0.410 1.310 0.490 1.790 ;
        RECT  0.170 1.310 0.410 3.380 ;
    END
END XNOR2XL

MACRO XNOR2X4
    CLASS CORE ;
    FOREIGN XNOR2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ XNOR2XL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  10.660 3.030 10.670 3.430 ;
        RECT  10.670 2.940 10.680 4.340 ;
        RECT  10.600 1.390 10.800 1.790 ;
        RECT  10.680 2.900 11.040 4.340 ;
        RECT  10.800 1.380 11.040 1.800 ;
        RECT  11.040 1.380 11.110 4.340 ;
        RECT  11.110 1.380 11.460 3.520 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.020 2.080 1.520 2.480 ;
        RECT  1.520 2.080 1.780 2.650 ;
        RECT  1.780 2.080 2.000 2.480 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.390 2.850 2.650 ;
        RECT  2.850 2.260 3.100 2.650 ;
        RECT  3.100 2.260 3.680 2.500 ;
        RECT  3.680 2.100 3.920 2.500 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.850 0.560 5.440 ;
        RECT  0.560 4.640 1.520 5.440 ;
        RECT  1.520 4.050 1.530 5.440 ;
        RECT  1.530 3.850 1.930 5.440 ;
        RECT  1.930 4.050 1.940 5.440 ;
        RECT  1.940 4.640 3.130 5.440 ;
        RECT  3.130 4.480 3.530 5.440 ;
        RECT  3.530 4.640 8.510 5.440 ;
        RECT  8.510 4.480 8.910 5.440 ;
        RECT  8.910 4.640 9.910 5.440 ;
        RECT  9.910 4.480 10.310 5.440 ;
        RECT  10.310 4.640 11.390 5.440 ;
        RECT  11.390 4.160 11.630 5.440 ;
        RECT  11.630 4.640 11.880 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.560 0.400 ;
        RECT  0.560 -0.400 0.570 0.840 ;
        RECT  0.570 -0.400 0.970 1.040 ;
        RECT  0.970 -0.400 0.980 0.840 ;
        RECT  0.980 -0.400 1.880 0.400 ;
        RECT  1.880 -0.400 1.890 0.840 ;
        RECT  1.890 -0.400 2.290 1.040 ;
        RECT  2.290 -0.400 2.300 0.840 ;
        RECT  2.300 -0.400 3.230 0.400 ;
        RECT  3.230 -0.400 3.630 0.560 ;
        RECT  3.630 -0.400 8.490 0.400 ;
        RECT  8.490 -0.400 8.890 0.560 ;
        RECT  8.890 -0.400 9.930 0.400 ;
        RECT  9.930 -0.400 10.330 0.560 ;
        RECT  10.330 -0.400 11.240 0.400 ;
        RECT  11.240 -0.400 11.250 0.790 ;
        RECT  11.250 -0.400 11.650 0.990 ;
        RECT  11.650 -0.400 11.660 0.790 ;
        RECT  11.660 -0.400 11.880 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.250 2.190 10.800 2.590 ;
        RECT  10.010 0.870 10.250 4.180 ;
        RECT  8.160 0.870 10.010 1.110 ;
        RECT  8.170 3.940 10.010 4.180 ;
        RECT  9.490 1.390 9.730 3.420 ;
        RECT  9.260 1.390 9.490 1.790 ;
        RECT  9.180 3.020 9.490 3.420 ;
        RECT  7.690 1.540 9.260 1.780 ;
        RECT  8.900 2.310 9.250 2.710 ;
        RECT  8.850 2.310 8.900 3.500 ;
        RECT  8.660 2.470 8.850 3.500 ;
        RECT  7.410 3.260 8.660 3.500 ;
        RECT  7.770 3.790 8.170 4.190 ;
        RECT  8.080 0.860 8.160 1.260 ;
        RECT  7.760 0.800 8.080 1.260 ;
        RECT  6.650 3.900 7.770 4.140 ;
        RECT  6.640 0.800 7.760 1.040 ;
        RECT  7.450 1.540 7.690 2.980 ;
        RECT  7.400 1.540 7.450 1.780 ;
        RECT  5.830 2.740 7.450 2.980 ;
        RECT  7.010 3.260 7.410 3.660 ;
        RECT  7.000 1.320 7.400 1.780 ;
        RECT  6.810 2.060 7.210 2.460 ;
        RECT  2.750 3.300 7.010 3.540 ;
        RECT  4.520 2.220 6.810 2.460 ;
        RECT  6.410 3.820 6.650 4.140 ;
        RECT  6.450 0.800 6.640 1.370 ;
        RECT  6.210 0.800 6.450 1.840 ;
        RECT  4.610 3.820 6.410 4.060 ;
        RECT  5.120 1.600 6.210 1.840 ;
        RECT  5.480 0.870 5.880 1.320 ;
        RECT  5.590 2.740 5.830 3.020 ;
        RECT  5.430 2.780 5.590 3.020 ;
        RECT  2.960 0.870 5.480 1.110 ;
        RECT  4.720 1.420 5.120 1.840 ;
        RECT  4.440 2.220 4.520 3.020 ;
        RECT  4.200 1.410 4.440 3.020 ;
        RECT  3.980 1.410 4.200 1.650 ;
        RECT  3.870 2.780 4.200 3.020 ;
        RECT  2.760 0.870 2.960 1.740 ;
        RECT  2.720 0.870 2.760 1.750 ;
        RECT  2.550 3.020 2.750 3.540 ;
        RECT  2.480 1.330 2.720 1.750 ;
        RECT  2.480 3.010 2.550 3.540 ;
        RECT  2.410 1.330 2.480 3.540 ;
        RECT  2.240 1.330 2.410 3.430 ;
        RECT  1.420 1.330 2.240 1.750 ;
        RECT  1.010 3.010 2.240 3.430 ;
        RECT  1.220 1.340 1.420 1.740 ;
        RECT  0.810 3.020 1.010 3.420 ;
    END
END XNOR2X4

MACRO XNOR2X2
    CLASS CORE ;
    FOREIGN XNOR2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ XNOR2XL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.650 2.820 6.810 3.800 ;
        RECT  6.690 0.660 6.810 1.640 ;
        RECT  6.810 0.660 7.050 3.800 ;
        RECT  7.050 3.510 7.060 3.770 ;
        RECT  7.050 0.660 7.090 1.960 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 0.870 3.210 ;
        RECT  0.870 2.580 0.890 3.210 ;
        RECT  0.890 2.580 1.240 3.220 ;
        RECT  1.240 2.580 1.820 2.820 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.690 1.900 1.090 2.300 ;
        RECT  1.090 1.900 2.100 2.140 ;
        RECT  2.100 1.900 2.180 2.640 ;
        RECT  2.180 1.900 2.340 2.650 ;
        RECT  2.340 2.160 2.440 2.650 ;
        RECT  2.440 2.160 2.690 2.580 ;
        RECT  2.690 2.170 2.810 2.570 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.960 5.440 ;
        RECT  0.960 4.480 1.360 5.440 ;
        RECT  1.360 4.640 2.490 5.440 ;
        RECT  2.490 3.930 2.890 5.440 ;
        RECT  2.890 4.640 5.830 5.440 ;
        RECT  5.830 4.480 6.230 5.440 ;
        RECT  6.230 4.640 7.260 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.830 0.400 ;
        RECT  0.830 -0.400 1.230 0.560 ;
        RECT  1.230 -0.400 2.470 0.400 ;
        RECT  2.470 -0.400 2.870 0.560 ;
        RECT  2.870 -0.400 5.870 0.400 ;
        RECT  5.870 -0.400 6.270 0.560 ;
        RECT  6.270 -0.400 7.260 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.890 1.980 6.570 2.220 ;
        RECT  5.650 0.860 5.890 2.220 ;
        RECT  5.570 2.620 5.810 4.120 ;
        RECT  4.810 0.860 5.650 1.100 ;
        RECT  5.380 3.880 5.570 4.120 ;
        RECT  5.140 3.880 5.380 4.370 ;
        RECT  5.330 1.380 5.370 1.780 ;
        RECT  5.090 1.380 5.330 3.590 ;
        RECT  3.610 4.130 5.140 4.370 ;
        RECT  4.570 0.860 4.810 3.850 ;
        RECT  4.290 1.050 4.570 1.450 ;
        RECT  3.930 3.610 4.570 3.850 ;
        RECT  4.050 2.010 4.290 3.330 ;
        RECT  3.850 2.010 4.050 2.250 ;
        RECT  3.610 3.090 4.050 3.330 ;
        RECT  3.610 0.860 3.850 2.250 ;
        RECT  3.330 2.540 3.810 2.780 ;
        RECT  2.050 0.860 3.610 1.100 ;
        RECT  3.330 3.090 3.610 4.370 ;
        RECT  3.090 1.380 3.330 2.780 ;
        RECT  3.210 3.240 3.330 4.140 ;
        RECT  2.050 3.350 3.210 3.590 ;
        RECT  0.570 1.380 3.090 1.620 ;
        RECT  1.650 0.790 2.050 1.100 ;
        RECT  1.650 3.190 2.050 3.590 ;
        RECT  0.390 1.220 0.570 1.620 ;
        RECT  0.390 3.240 0.480 3.640 ;
        RECT  0.150 1.220 0.390 3.640 ;
    END
END XNOR2X2

MACRO XNOR2X1
    CLASS CORE ;
    FOREIGN XNOR2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ XNOR2XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.820 2.950 5.040 3.210 ;
        RECT  5.040 2.950 5.450 3.490 ;
        RECT  5.450 1.200 5.610 3.490 ;
        RECT  5.610 1.200 5.690 3.190 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 1.980 1.870 2.660 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 1.750 1.120 2.170 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.610 5.440 ;
        RECT  0.610 4.020 0.620 5.440 ;
        RECT  0.620 3.900 1.020 5.440 ;
        RECT  1.020 4.020 1.030 5.440 ;
        RECT  1.030 4.640 4.220 5.440 ;
        RECT  4.220 4.480 4.620 5.440 ;
        RECT  4.620 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.340 0.400 ;
        RECT  0.340 -0.400 0.740 0.560 ;
        RECT  0.740 -0.400 4.570 0.400 ;
        RECT  4.570 -0.400 4.970 0.560 ;
        RECT  4.970 -0.400 5.940 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.850 0.860 5.090 2.570 ;
        RECT  3.510 0.860 4.850 1.100 ;
        RECT  3.790 1.380 4.030 3.150 ;
        RECT  3.700 3.740 3.980 3.980 ;
        RECT  3.340 2.910 3.790 3.150 ;
        RECT  3.460 3.510 3.700 3.980 ;
        RECT  3.270 0.860 3.510 1.430 ;
        RECT  2.380 3.510 3.460 3.750 ;
        RECT  2.900 1.190 3.270 1.430 ;
        RECT  1.280 0.670 2.990 0.910 ;
        RECT  2.660 1.190 2.900 3.230 ;
        RECT  1.540 4.030 2.660 4.270 ;
        RECT  2.140 1.440 2.380 3.750 ;
        RECT  1.970 1.440 2.140 1.680 ;
        RECT  1.820 3.010 2.140 3.410 ;
        RECT  1.570 1.220 1.970 1.680 ;
        RECT  1.300 3.140 1.540 4.270 ;
        RECT  0.570 3.140 1.300 3.380 ;
        RECT  1.040 0.670 1.280 1.100 ;
        RECT  0.490 0.860 1.040 1.100 ;
        RECT  0.410 2.980 0.570 3.380 ;
        RECT  0.410 0.860 0.490 1.400 ;
        RECT  0.200 0.860 0.410 3.380 ;
        RECT  0.170 1.160 0.200 3.380 ;
    END
END XNOR2X1

MACRO TTLATXL
    CLASS CORE ;
    FOREIGN TTLATXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.240 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  6.140 2.950 6.150 3.210 ;
        RECT  6.150 1.380 6.160 3.330 ;
        RECT  6.160 1.380 6.390 3.340 ;
        RECT  6.390 2.940 6.560 3.340 ;
        RECT  6.390 1.380 6.620 1.780 ;
        END
    END Q
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.710 2.060 7.150 2.660 ;
        END
    END OE
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  8.030 2.240 8.460 2.660 ;
        RECT  8.460 2.250 8.550 2.650 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.940 2.360 2.530 2.760 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.720 5.440 ;
        RECT  1.720 4.480 2.120 5.440 ;
        RECT  2.120 4.640 4.750 5.440 ;
        RECT  4.540 3.400 4.750 3.800 ;
        RECT  4.750 3.400 4.780 5.440 ;
        RECT  4.780 3.420 5.110 5.440 ;
        RECT  5.110 4.640 7.790 5.440 ;
        RECT  7.790 3.450 8.190 5.440 ;
        RECT  8.190 4.640 9.240 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.370 0.400 ;
        RECT  0.370 -0.400 1.910 0.560 ;
        RECT  1.910 -0.400 4.510 0.400 ;
        RECT  4.510 -0.400 4.910 0.560 ;
        RECT  4.910 -0.400 7.780 0.400 ;
        RECT  7.780 -0.400 8.180 0.560 ;
        RECT  8.180 -0.400 9.240 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  8.910 1.400 9.070 3.320 ;
        RECT  8.830 0.860 8.910 3.320 ;
        RECT  8.670 0.860 8.830 1.800 ;
        RECT  8.670 2.920 8.830 3.320 ;
        RECT  4.190 0.860 8.670 1.100 ;
        RECT  7.420 1.560 7.660 3.160 ;
        RECT  7.360 1.560 7.420 1.800 ;
        RECT  7.300 2.920 7.420 3.160 ;
        RECT  6.960 1.400 7.360 1.800 ;
        RECT  7.140 2.920 7.300 3.320 ;
        RECT  6.900 2.920 7.140 3.850 ;
        RECT  6.250 3.610 6.900 3.850 ;
        RECT  5.850 3.610 6.250 4.010 ;
        RECT  5.500 1.380 5.740 3.150 ;
        RECT  5.340 1.380 5.500 1.780 ;
        RECT  5.280 2.750 5.500 3.150 ;
        RECT  4.820 2.070 5.220 2.470 ;
        RECT  4.240 2.150 4.820 2.390 ;
        RECT  2.640 4.080 4.470 4.320 ;
        RECT  4.000 1.590 4.240 3.800 ;
        RECT  3.950 0.670 4.190 1.100 ;
        RECT  3.670 1.590 4.000 1.830 ;
        RECT  3.160 3.560 4.000 3.800 ;
        RECT  2.640 0.670 3.950 0.910 ;
        RECT  3.460 2.880 3.700 3.280 ;
        RECT  3.430 1.190 3.670 1.830 ;
        RECT  3.130 2.880 3.460 3.120 ;
        RECT  3.050 1.190 3.430 1.430 ;
        RECT  2.920 3.420 3.160 3.800 ;
        RECT  2.890 1.720 3.130 3.120 ;
        RECT  0.920 3.420 2.920 3.660 ;
        RECT  1.500 1.720 2.890 1.960 ;
        RECT  2.400 0.670 2.640 1.150 ;
        RECT  2.400 3.940 2.640 4.320 ;
        RECT  1.400 0.910 2.400 1.150 ;
        RECT  1.440 3.940 2.400 4.180 ;
        RECT  1.290 1.470 1.500 1.960 ;
        RECT  1.200 3.940 1.440 4.360 ;
        RECT  1.050 1.470 1.290 3.100 ;
        RECT  0.400 4.120 1.200 4.360 ;
        RECT  0.770 2.860 1.050 3.100 ;
        RECT  0.680 3.420 0.920 3.850 ;
        RECT  0.400 1.390 0.620 1.790 ;
        RECT  0.160 1.390 0.400 4.360 ;
    END
END TTLATXL

MACRO TTLATX4
    CLASS CORE ;
    FOREIGN TTLATX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TTLATXL ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  10.630 3.130 10.890 3.530 ;
        RECT  10.890 2.840 11.330 3.780 ;
        RECT  11.330 2.380 12.100 3.780 ;
        RECT  10.600 1.200 12.100 1.440 ;
        RECT  12.100 1.200 12.210 3.780 ;
        RECT  12.210 1.200 12.340 3.530 ;
        RECT  12.340 1.390 12.540 1.790 ;
        RECT  12.340 3.130 12.550 3.530 ;
        END
    END Q
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  13.400 2.950 13.410 3.210 ;
        RECT  13.410 2.230 13.650 3.210 ;
        RECT  13.650 2.950 13.660 3.210 ;
        END
    END OE
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  14.060 1.830 14.070 2.090 ;
        RECT  14.070 1.830 14.320 2.310 ;
        RECT  14.320 2.070 14.770 2.310 ;
        RECT  14.770 2.070 15.010 2.470 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.790 1.920 3.950 2.320 ;
        RECT  3.950 1.850 4.160 2.320 ;
        RECT  4.160 1.830 4.190 2.320 ;
        RECT  4.190 1.830 4.420 2.090 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.040 5.440 ;
        RECT  1.040 4.480 1.440 5.440 ;
        RECT  1.440 4.640 3.600 5.440 ;
        RECT  3.600 4.480 4.000 5.440 ;
        RECT  4.000 4.640 5.400 5.440 ;
        RECT  5.400 4.480 5.800 5.440 ;
        RECT  5.800 4.640 7.480 5.440 ;
        RECT  7.480 4.010 7.880 5.440 ;
        RECT  7.880 4.640 9.140 5.440 ;
        RECT  9.140 4.010 9.540 5.440 ;
        RECT  9.540 4.640 14.490 5.440 ;
        RECT  14.490 3.060 14.890 5.440 ;
        RECT  14.890 4.640 15.840 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.290 0.400 ;
        RECT  0.290 -0.400 0.690 0.560 ;
        RECT  0.690 -0.400 1.890 0.400 ;
        RECT  1.890 -0.400 2.290 0.560 ;
        RECT  2.290 -0.400 6.360 0.400 ;
        RECT  6.360 -0.400 6.760 0.560 ;
        RECT  6.760 -0.400 7.770 0.400 ;
        RECT  7.770 -0.400 8.170 0.560 ;
        RECT  8.170 -0.400 9.170 0.400 ;
        RECT  9.170 -0.400 9.570 0.560 ;
        RECT  9.570 -0.400 13.980 0.400 ;
        RECT  13.980 -0.400 14.380 0.560 ;
        RECT  14.380 -0.400 15.840 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  15.530 2.740 15.650 4.140 ;
        RECT  15.290 1.550 15.530 4.140 ;
        RECT  15.120 1.550 15.290 1.790 ;
        RECT  15.250 2.740 15.290 4.140 ;
        RECT  14.880 0.750 15.120 1.790 ;
        RECT  13.490 0.870 14.880 1.110 ;
        RECT  13.730 3.490 14.130 3.890 ;
        RECT  13.060 3.490 13.730 3.730 ;
        RECT  13.250 0.680 13.490 1.110 ;
        RECT  13.070 1.400 13.470 1.800 ;
        RECT  10.290 4.050 13.260 4.290 ;
        RECT  10.160 0.680 13.250 0.920 ;
        RECT  13.060 1.560 13.070 1.800 ;
        RECT  12.820 1.560 13.060 3.730 ;
        RECT  12.800 2.440 12.820 3.730 ;
        RECT  12.690 2.440 12.800 2.840 ;
        RECT  10.260 1.720 11.820 1.960 ;
        RECT  10.260 3.120 10.290 4.290 ;
        RECT  10.240 1.720 10.260 4.290 ;
        RECT  10.050 1.390 10.240 4.290 ;
        RECT  9.920 0.680 10.160 1.100 ;
        RECT  9.890 1.390 10.050 3.520 ;
        RECT  5.970 0.860 9.920 1.100 ;
        RECT  9.840 1.390 9.890 3.180 ;
        RECT  8.840 1.470 9.840 1.710 ;
        RECT  6.980 2.780 9.840 3.180 ;
        RECT  6.880 2.100 9.150 2.500 ;
        RECT  8.440 1.390 8.840 1.790 ;
        RECT  7.500 1.470 8.440 1.710 ;
        RECT  7.100 1.390 7.500 1.790 ;
        RECT  6.740 2.080 6.880 2.500 ;
        RECT  6.670 3.890 6.760 4.130 ;
        RECT  6.630 2.080 6.740 3.530 ;
        RECT  6.360 3.890 6.670 4.180 ;
        RECT  6.500 1.380 6.630 3.530 ;
        RECT  6.390 1.380 6.500 2.320 ;
        RECT  5.490 3.290 6.500 3.530 ;
        RECT  5.450 1.380 6.390 1.620 ;
        RECT  0.480 3.940 6.360 4.180 ;
        RECT  6.020 2.600 6.260 3.010 ;
        RECT  5.050 2.600 6.020 2.840 ;
        RECT  5.730 0.760 5.970 1.100 ;
        RECT  2.810 0.760 5.730 1.000 ;
        RECT  5.250 3.120 5.490 3.530 ;
        RECT  5.090 1.330 5.450 1.620 ;
        RECT  5.070 3.120 5.250 3.500 ;
        RECT  4.850 1.310 5.090 1.620 ;
        RECT  2.750 3.260 5.070 3.500 ;
        RECT  4.810 1.870 5.050 2.840 ;
        RECT  3.410 1.310 4.850 1.550 ;
        RECT  3.160 2.600 4.810 2.840 ;
        RECT  3.170 1.310 3.410 1.620 ;
        RECT  2.500 1.380 3.170 1.620 ;
        RECT  2.920 1.950 3.160 2.840 ;
        RECT  2.760 1.950 2.920 2.280 ;
        RECT  2.570 0.760 2.810 1.100 ;
        RECT  1.950 2.040 2.760 2.280 ;
        RECT  2.350 3.260 2.750 3.660 ;
        RECT  2.220 0.860 2.570 1.100 ;
        RECT  1.020 3.420 2.350 3.660 ;
        RECT  1.980 0.860 2.220 1.760 ;
        RECT  1.950 2.820 2.030 3.060 ;
        RECT  1.820 1.520 1.980 1.760 ;
        RECT  1.710 2.040 1.950 3.060 ;
        RECT  1.540 2.040 1.710 2.280 ;
        RECT  1.630 2.820 1.710 3.060 ;
        RECT  1.300 0.950 1.540 2.280 ;
        RECT  1.070 0.950 1.300 1.190 ;
        RECT  0.990 2.260 1.020 3.660 ;
        RECT  0.780 2.180 0.990 3.660 ;
        RECT  0.750 2.180 0.780 2.580 ;
        RECT  0.480 1.390 0.620 1.790 ;
        RECT  0.240 1.390 0.480 4.180 ;
        RECT  0.220 1.390 0.240 1.790 ;
    END
END TTLATX4

MACRO TTLATX2
    CLASS CORE ;
    FOREIGN TTLATX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TTLATXL ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  8.780 2.950 8.830 3.210 ;
        RECT  8.830 2.640 8.930 3.210 ;
        RECT  8.930 1.380 9.040 3.210 ;
        RECT  9.040 1.380 9.170 3.200 ;
        RECT  9.170 1.380 9.330 1.780 ;
        END
    END Q
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  10.580 2.420 10.670 2.820 ;
        RECT  10.670 2.420 10.740 2.940 ;
        RECT  10.740 2.420 10.760 3.190 ;
        RECT  10.760 2.420 10.980 3.210 ;
        RECT  10.980 2.950 11.020 3.210 ;
        END
    END OE
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  11.360 2.070 11.420 2.470 ;
        RECT  11.420 1.830 11.680 2.470 ;
        RECT  11.680 2.070 11.760 2.470 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.710 1.830 4.110 2.320 ;
        RECT  4.110 1.830 4.420 2.090 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.750 5.440 ;
        RECT  1.750 4.480 2.150 5.440 ;
        RECT  2.150 4.640 3.490 5.440 ;
        RECT  3.490 4.100 3.890 5.440 ;
        RECT  3.890 4.640 5.220 5.440 ;
        RECT  5.220 4.480 5.620 5.440 ;
        RECT  5.620 4.640 7.340 5.440 ;
        RECT  7.340 4.010 7.740 5.440 ;
        RECT  7.740 4.640 11.090 5.440 ;
        RECT  11.090 3.500 11.490 5.440 ;
        RECT  11.490 4.640 12.540 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.200 0.400 ;
        RECT  0.200 -0.400 2.300 0.560 ;
        RECT  2.300 -0.400 6.170 0.400 ;
        RECT  6.170 -0.400 6.570 0.560 ;
        RECT  6.570 -0.400 7.500 0.400 ;
        RECT  7.500 -0.400 7.900 0.560 ;
        RECT  7.900 -0.400 11.210 0.400 ;
        RECT  11.210 -0.400 11.610 0.560 ;
        RECT  11.610 -0.400 12.540 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.210 0.860 12.290 3.450 ;
        RECT  12.050 0.860 12.210 3.780 ;
        RECT  5.890 0.860 12.050 1.100 ;
        RECT  11.810 2.880 12.050 3.780 ;
        RECT  10.670 1.400 10.830 1.800 ;
        RECT  10.420 3.490 10.760 3.730 ;
        RECT  10.430 1.400 10.670 2.140 ;
        RECT  10.420 4.060 10.580 4.300 ;
        RECT  10.290 1.900 10.430 2.140 ;
        RECT  10.290 3.450 10.420 4.300 ;
        RECT  10.180 1.900 10.290 4.300 ;
        RECT  10.050 1.900 10.180 3.690 ;
        RECT  9.810 1.380 10.090 1.620 ;
        RECT  9.810 3.930 9.940 4.330 ;
        RECT  9.700 1.380 9.810 4.330 ;
        RECT  9.570 1.380 9.700 4.250 ;
        RECT  8.500 3.490 9.570 3.730 ;
        RECT  8.420 1.390 8.570 1.790 ;
        RECT  8.420 3.490 8.500 3.900 ;
        RECT  8.180 1.390 8.420 3.900 ;
        RECT  8.170 1.390 8.180 1.790 ;
        RECT  8.100 2.780 8.180 3.900 ;
        RECT  7.230 1.480 8.170 1.720 ;
        RECT  7.050 2.780 8.100 3.020 ;
        RECT  6.570 2.080 7.900 2.500 ;
        RECT  6.830 1.400 7.230 1.800 ;
        RECT  6.810 2.780 7.050 3.180 ;
        RECT  6.510 3.850 6.590 4.090 ;
        RECT  6.330 1.380 6.570 3.530 ;
        RECT  6.420 3.850 6.510 4.120 ;
        RECT  6.180 3.850 6.420 4.180 ;
        RECT  5.370 1.380 6.330 1.620 ;
        RECT  5.470 3.290 6.330 3.530 ;
        RECT  4.390 3.940 6.180 4.180 ;
        RECT  5.850 2.600 6.090 3.010 ;
        RECT  5.650 0.670 5.890 1.100 ;
        RECT  4.990 2.600 5.850 2.840 ;
        RECT  2.810 0.670 5.650 0.910 ;
        RECT  5.230 3.090 5.470 3.530 ;
        RECT  5.030 1.330 5.370 1.620 ;
        RECT  2.690 3.090 5.230 3.330 ;
        RECT  4.790 1.190 5.030 1.620 ;
        RECT  4.750 1.870 4.990 2.840 ;
        RECT  3.330 1.190 4.790 1.430 ;
        RECT  3.050 2.600 4.750 2.840 ;
        RECT  4.150 3.600 4.390 4.180 ;
        RECT  3.180 3.600 4.150 3.840 ;
        RECT  3.090 1.190 3.330 1.630 ;
        RECT  2.940 3.600 3.180 4.180 ;
        RECT  2.420 1.390 3.090 1.630 ;
        RECT  3.050 1.950 3.080 2.190 ;
        RECT  2.810 1.950 3.050 2.840 ;
        RECT  1.470 3.940 2.940 4.180 ;
        RECT  2.570 0.670 2.810 1.100 ;
        RECT  1.490 1.950 2.810 2.190 ;
        RECT  2.540 3.080 2.690 3.480 ;
        RECT  1.720 0.860 2.570 1.100 ;
        RECT  2.290 3.080 2.540 3.660 ;
        RECT  0.940 3.420 2.290 3.660 ;
        RECT  1.310 0.860 1.720 1.150 ;
        RECT  1.470 1.480 1.490 2.190 ;
        RECT  1.230 1.480 1.470 3.090 ;
        RECT  1.230 3.940 1.470 4.360 ;
        RECT  1.090 1.480 1.230 1.720 ;
        RECT  0.950 2.850 1.230 3.090 ;
        RECT  0.420 4.120 1.230 4.360 ;
        RECT  0.700 3.420 0.940 3.860 ;
        RECT  0.420 1.390 0.620 1.790 ;
        RECT  0.180 1.390 0.420 4.360 ;
    END
END TTLATX2

MACRO TTLATX1
    CLASS CORE ;
    FOREIGN TTLATX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TTLATXL ;
    SIZE 9.240 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Q
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  5.480 3.510 5.590 3.770 ;
        RECT  5.590 3.500 5.950 3.780 ;
        RECT  5.950 3.500 6.100 4.290 ;
        RECT  6.100 1.380 6.340 4.290 ;
        RECT  6.340 3.890 6.350 4.290 ;
        RECT  6.340 1.380 6.500 1.780 ;
        END
    END Q
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.710 2.060 7.150 2.660 ;
        END
    END OE
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  8.030 2.240 8.460 2.660 ;
        RECT  8.460 2.250 8.550 2.650 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.090 2.360 2.490 2.980 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.720 5.440 ;
        RECT  1.720 4.480 2.120 5.440 ;
        RECT  2.120 4.640 4.740 5.440 ;
        RECT  4.740 3.900 4.750 5.440 ;
        RECT  4.750 3.890 5.120 5.440 ;
        RECT  5.120 4.640 7.930 5.440 ;
        RECT  7.930 2.920 8.350 5.440 ;
        RECT  8.350 4.640 9.240 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.380 0.400 ;
        RECT  0.380 -0.400 2.140 0.560 ;
        RECT  2.140 -0.400 4.510 0.400 ;
        RECT  4.510 -0.400 4.910 0.560 ;
        RECT  4.910 -0.400 7.770 0.400 ;
        RECT  7.770 -0.400 8.170 0.560 ;
        RECT  8.170 -0.400 9.240 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  8.910 1.350 9.070 3.330 ;
        RECT  8.830 0.860 8.910 3.330 ;
        RECT  8.670 0.860 8.830 1.800 ;
        RECT  8.670 2.930 8.830 3.330 ;
        RECT  4.190 0.860 8.670 1.100 ;
        RECT  7.420 1.560 7.660 3.160 ;
        RECT  7.260 1.560 7.420 1.800 ;
        RECT  7.410 2.920 7.420 3.160 ;
        RECT  7.250 2.920 7.410 3.320 ;
        RECT  6.860 1.400 7.260 1.800 ;
        RECT  7.020 2.920 7.250 4.200 ;
        RECT  7.010 2.920 7.020 4.360 ;
        RECT  6.620 3.960 7.010 4.360 ;
        RECT  5.500 1.380 5.740 3.180 ;
        RECT  5.340 1.380 5.500 1.780 ;
        RECT  5.280 2.780 5.500 3.180 ;
        RECT  4.820 2.090 5.220 2.490 ;
        RECT  4.240 2.170 4.820 2.410 ;
        RECT  2.640 4.080 4.470 4.320 ;
        RECT  4.000 1.590 4.240 3.800 ;
        RECT  3.950 0.670 4.190 1.100 ;
        RECT  3.670 1.590 4.000 1.830 ;
        RECT  3.160 3.560 4.000 3.800 ;
        RECT  2.640 0.670 3.950 0.910 ;
        RECT  3.460 2.880 3.700 3.280 ;
        RECT  3.430 1.190 3.670 1.830 ;
        RECT  3.130 2.880 3.460 3.120 ;
        RECT  3.050 1.190 3.430 1.430 ;
        RECT  2.920 3.420 3.160 3.800 ;
        RECT  2.890 1.700 3.130 3.120 ;
        RECT  0.920 3.420 2.920 3.660 ;
        RECT  1.490 1.700 2.890 1.940 ;
        RECT  2.400 0.670 2.640 1.150 ;
        RECT  2.400 3.940 2.640 4.320 ;
        RECT  1.390 0.910 2.400 1.150 ;
        RECT  1.440 3.940 2.400 4.180 ;
        RECT  1.290 1.470 1.490 1.940 ;
        RECT  1.200 3.940 1.440 4.360 ;
        RECT  1.050 1.470 1.290 3.100 ;
        RECT  0.400 4.120 1.200 4.360 ;
        RECT  0.770 2.860 1.050 3.100 ;
        RECT  0.680 3.420 0.920 3.850 ;
        RECT  0.400 1.390 0.620 1.790 ;
        RECT  0.160 1.390 0.400 4.360 ;
    END
END TTLATX1

MACRO TLATSRXL
    CLASS CORE ;
    FOREIGN TLATSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.180 1.830 0.600 2.600 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.460 1.820 3.860 2.410 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  10.650 2.990 10.770 3.390 ;
        RECT  10.760 2.390 10.770 2.650 ;
        RECT  10.650 1.240 10.770 1.820 ;
        RECT  10.770 1.240 11.010 3.390 ;
        RECT  11.010 2.390 11.020 2.650 ;
        RECT  11.010 2.990 11.050 3.390 ;
        RECT  11.010 1.240 11.050 1.960 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.250 2.950 9.560 3.350 ;
        RECT  9.250 1.470 9.560 1.710 ;
        RECT  9.560 1.470 9.800 3.350 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  6.140 1.830 6.150 2.090 ;
        RECT  6.150 1.830 6.400 2.230 ;
        RECT  6.400 1.990 6.520 2.230 ;
        RECT  6.520 1.990 6.920 2.390 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.740 1.990 2.840 2.390 ;
        RECT  2.840 1.990 3.100 2.650 ;
        RECT  3.100 1.990 3.140 2.520 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.790 0.560 5.440 ;
        RECT  0.560 4.640 3.100 5.440 ;
        RECT  3.100 4.060 3.500 5.440 ;
        RECT  3.500 4.640 6.500 5.440 ;
        RECT  6.500 4.480 6.900 5.440 ;
        RECT  6.900 4.640 8.410 5.440 ;
        RECT  8.410 4.480 8.810 5.440 ;
        RECT  8.810 4.640 10.040 5.440 ;
        RECT  10.040 4.480 10.440 5.440 ;
        RECT  10.440 4.640 11.220 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 2.450 0.400 ;
        RECT  2.450 -0.400 2.850 0.560 ;
        RECT  2.850 -0.400 6.170 0.400 ;
        RECT  6.170 -0.400 6.570 0.560 ;
        RECT  6.570 -0.400 8.450 0.400 ;
        RECT  8.450 -0.400 8.690 1.860 ;
        RECT  8.690 -0.400 9.980 0.400 ;
        RECT  9.980 -0.400 10.380 0.560 ;
        RECT  10.380 -0.400 11.220 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.110 0.880 10.350 4.020 ;
        RECT  9.650 0.880 10.110 1.120 ;
        RECT  9.710 3.780 10.110 4.020 ;
        RECT  9.470 3.780 9.710 4.370 ;
        RECT  9.250 0.720 9.650 1.120 ;
        RECT  9.310 3.940 9.470 4.370 ;
        RECT  6.210 3.940 9.310 4.180 ;
        RECT  8.930 2.210 9.230 2.610 ;
        RECT  8.830 2.210 8.930 3.660 ;
        RECT  8.690 2.220 8.830 3.660 ;
        RECT  4.710 3.420 8.690 3.660 ;
        RECT  7.930 0.680 8.170 3.140 ;
        RECT  7.710 0.680 7.930 1.100 ;
        RECT  7.770 2.900 7.930 3.140 ;
        RECT  5.590 0.860 7.710 1.100 ;
        RECT  7.470 2.020 7.650 2.420 ;
        RECT  7.230 1.420 7.470 3.140 ;
        RECT  7.000 1.420 7.230 1.660 ;
        RECT  4.620 2.900 7.230 3.140 ;
        RECT  5.810 3.940 6.210 4.350 ;
        RECT  5.350 0.860 5.590 2.620 ;
        RECT  4.900 2.380 5.350 2.620 ;
        RECT  4.620 1.580 5.070 1.980 ;
        RECT  4.410 0.860 4.810 1.250 ;
        RECT  4.390 3.420 4.710 3.780 ;
        RECT  4.360 1.580 4.620 3.140 ;
        RECT  2.800 0.860 4.410 1.100 ;
        RECT  1.890 3.540 4.390 3.780 ;
        RECT  4.090 2.900 4.360 3.140 ;
        RECT  3.850 2.900 4.090 3.260 ;
        RECT  2.410 3.020 3.850 3.260 ;
        RECT  2.560 0.860 2.800 1.560 ;
        RECT  1.670 1.320 2.560 1.560 ;
        RECT  2.170 2.040 2.410 3.260 ;
        RECT  1.950 2.040 2.170 2.440 ;
        RECT  1.150 0.770 2.160 1.010 ;
        RECT  1.670 3.090 1.890 3.780 ;
        RECT  1.150 4.060 1.770 4.300 ;
        RECT  1.650 1.320 1.670 3.780 ;
        RECT  1.430 1.320 1.650 3.330 ;
        RECT  0.910 0.770 1.150 4.300 ;
    END
END TLATSRXL

MACRO TLATSRX4
    CLASS CORE ;
    FOREIGN TLATSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATSRXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.520 1.780 1.120 2.200 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.780 1.830 8.790 2.090 ;
        RECT  8.790 1.830 9.040 2.420 ;
        RECT  9.040 1.840 9.110 2.420 ;
        RECT  9.110 2.020 9.190 2.420 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.290 1.820 15.330 3.220 ;
        RECT  15.330 1.220 15.640 3.220 ;
        RECT  15.640 1.220 15.730 3.250 ;
        RECT  15.730 2.850 16.040 3.250 ;
        RECT  15.730 1.220 16.040 1.630 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.970 1.820 14.100 3.220 ;
        RECT  14.100 1.230 14.420 3.250 ;
        RECT  14.420 2.850 14.500 3.250 ;
        RECT  14.420 1.230 14.500 1.630 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  10.010 2.100 10.100 2.500 ;
        RECT  10.100 1.830 10.360 2.500 ;
        RECT  10.360 2.100 10.410 2.500 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.510 2.090 ;
        RECT  3.510 1.830 3.750 2.620 ;
        RECT  3.750 1.830 3.760 2.090 ;
        RECT  3.750 2.380 5.270 2.620 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.930 5.440 ;
        RECT  0.930 3.200 1.330 5.440 ;
        RECT  1.330 4.640 6.350 5.440 ;
        RECT  6.350 4.480 6.750 5.440 ;
        RECT  6.750 4.640 10.010 5.440 ;
        RECT  10.010 4.480 10.410 5.440 ;
        RECT  10.410 4.640 11.890 5.440 ;
        RECT  11.890 4.480 12.290 5.440 ;
        RECT  12.290 4.640 13.360 5.440 ;
        RECT  13.360 4.480 13.760 5.440 ;
        RECT  13.760 4.640 14.890 5.440 ;
        RECT  14.890 4.210 15.290 5.440 ;
        RECT  15.290 4.640 16.310 5.440 ;
        RECT  16.310 4.210 16.710 5.440 ;
        RECT  16.710 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.200 0.400 ;
        RECT  1.200 -0.400 1.600 0.560 ;
        RECT  1.600 -0.400 2.960 0.400 ;
        RECT  2.960 -0.400 3.360 0.560 ;
        RECT  3.360 -0.400 5.850 0.400 ;
        RECT  5.850 -0.400 6.250 0.870 ;
        RECT  6.250 -0.400 9.130 0.400 ;
        RECT  9.130 -0.400 9.530 0.560 ;
        RECT  9.530 -0.400 12.050 0.400 ;
        RECT  12.050 -0.400 12.450 0.560 ;
        RECT  12.450 -0.400 13.490 0.400 ;
        RECT  13.490 -0.400 13.890 0.950 ;
        RECT  13.890 -0.400 14.920 0.400 ;
        RECT  14.920 -0.400 15.320 0.950 ;
        RECT  15.320 -0.400 16.310 0.400 ;
        RECT  16.310 -0.400 16.710 0.950 ;
        RECT  16.710 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.320 2.170 16.560 3.860 ;
        RECT  13.020 3.620 16.320 3.860 ;
        RECT  13.300 1.390 13.540 3.040 ;
        RECT  13.060 1.390 13.300 1.630 ;
        RECT  13.020 2.800 13.300 3.040 ;
        RECT  12.660 1.230 13.060 1.630 ;
        RECT  12.780 2.800 13.020 4.180 ;
        RECT  12.590 2.120 12.990 2.520 ;
        RECT  9.710 3.940 12.780 4.180 ;
        RECT  12.480 2.280 12.590 2.520 ;
        RECT  12.240 2.280 12.480 3.660 ;
        RECT  2.550 3.420 12.240 3.660 ;
        RECT  11.680 0.860 11.920 3.140 ;
        RECT  11.490 0.860 11.680 1.100 ;
        RECT  11.280 2.900 11.680 3.140 ;
        RECT  11.240 0.670 11.490 1.100 ;
        RECT  11.000 1.680 11.360 2.080 ;
        RECT  10.050 0.670 11.240 0.910 ;
        RECT  10.760 1.190 11.000 3.140 ;
        RECT  10.330 1.190 10.760 1.430 ;
        RECT  8.390 2.900 10.760 3.140 ;
        RECT  9.810 0.670 10.050 1.430 ;
        RECT  7.790 1.190 9.810 1.430 ;
        RECT  9.390 3.940 9.710 4.230 ;
        RECT  9.310 3.990 9.390 4.230 ;
        RECT  7.430 4.130 8.990 4.370 ;
        RECT  8.150 1.760 8.390 3.140 ;
        RECT  3.080 2.900 8.150 3.140 ;
        RECT  6.950 0.670 8.050 0.910 ;
        RECT  7.550 1.190 7.790 2.360 ;
        RECT  7.340 1.840 7.550 2.360 ;
        RECT  7.190 3.940 7.430 4.370 ;
        RECT  4.550 1.840 7.340 2.080 ;
        RECT  6.040 3.940 7.190 4.180 ;
        RECT  6.710 0.670 6.950 1.390 ;
        RECT  5.530 1.150 6.710 1.390 ;
        RECT  5.800 3.940 6.040 4.360 ;
        RECT  1.870 4.120 5.800 4.360 ;
        RECT  5.290 1.040 5.530 1.390 ;
        RECT  2.550 1.040 5.290 1.280 ;
        RECT  4.150 1.700 4.550 2.100 ;
        RECT  2.840 2.180 3.080 3.140 ;
        RECT  2.310 1.040 2.550 3.660 ;
        RECT  2.150 1.040 2.310 1.450 ;
        RECT  1.870 1.780 2.030 2.180 ;
        RECT  1.630 1.200 1.870 4.360 ;
        RECT  0.630 1.200 1.630 1.440 ;
        RECT  0.570 2.620 1.630 2.860 ;
        RECT  0.230 1.040 0.630 1.440 ;
        RECT  0.250 2.620 0.570 4.230 ;
        RECT  0.170 2.830 0.250 4.230 ;
    END
END TLATSRX4

MACRO TLATSRX2
    CLASS CORE ;
    FOREIGN TLATSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATSRXL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.190 1.900 0.200 2.420 ;
        RECT  0.200 1.830 0.460 2.420 ;
        RECT  0.460 1.900 0.590 2.420 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.510 2.070 3.670 2.470 ;
        RECT  3.670 1.860 3.910 2.470 ;
        RECT  3.910 1.860 4.160 2.100 ;
        RECT  4.160 1.830 4.400 2.100 ;
        RECT  4.400 1.830 4.420 2.090 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.340 1.260 11.390 3.390 ;
        RECT  11.390 1.180 11.630 3.390 ;
        RECT  11.630 1.460 11.640 3.020 ;
        RECT  11.640 2.390 11.680 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.440 2.950 9.700 3.210 ;
        RECT  9.700 2.960 10.070 3.200 ;
        RECT  10.070 2.880 10.300 3.280 ;
        RECT  9.700 1.410 10.300 1.650 ;
        RECT  10.300 1.410 10.470 3.280 ;
        RECT  10.470 1.410 10.540 3.120 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  6.140 1.830 6.160 2.090 ;
        RECT  6.160 1.830 6.400 2.610 ;
        RECT  6.400 2.370 6.950 2.610 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.790 1.530 2.840 1.930 ;
        RECT  2.840 1.530 3.100 2.090 ;
        RECT  3.100 1.530 3.110 2.080 ;
        RECT  3.110 1.530 3.190 1.930 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 3.250 5.440 ;
        RECT  3.250 3.790 3.650 5.440 ;
        RECT  3.650 4.640 6.570 5.440 ;
        RECT  6.570 4.480 6.970 5.440 ;
        RECT  6.970 4.640 8.470 5.440 ;
        RECT  8.470 4.480 8.870 5.440 ;
        RECT  8.870 4.640 10.700 5.440 ;
        RECT  10.700 4.190 11.100 5.440 ;
        RECT  11.100 4.640 11.880 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 2.460 0.400 ;
        RECT  2.460 -0.400 2.860 0.560 ;
        RECT  2.860 -0.400 6.350 0.400 ;
        RECT  6.350 -0.400 6.750 0.560 ;
        RECT  6.750 -0.400 8.370 0.400 ;
        RECT  8.370 -0.400 8.770 0.560 ;
        RECT  8.770 -0.400 10.590 0.400 ;
        RECT  10.590 -0.400 10.990 0.560 ;
        RECT  10.990 -0.400 11.880 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.820 0.880 11.060 3.860 ;
        RECT  10.110 0.880 10.820 1.120 ;
        RECT  9.750 3.620 10.820 3.860 ;
        RECT  9.870 0.670 10.110 1.120 ;
        RECT  9.060 2.040 10.030 2.440 ;
        RECT  9.140 0.670 9.870 0.910 ;
        RECT  9.340 3.620 9.750 4.180 ;
        RECT  6.290 3.940 9.340 4.180 ;
        RECT  8.910 2.040 9.060 3.660 ;
        RECT  8.820 2.200 8.910 3.660 ;
        RECT  4.390 3.420 8.820 3.660 ;
        RECT  8.300 0.860 8.540 3.140 ;
        RECT  8.020 0.860 8.300 1.100 ;
        RECT  7.860 2.900 8.300 3.140 ;
        RECT  7.620 0.670 8.020 1.100 ;
        RECT  7.490 1.900 8.020 2.300 ;
        RECT  5.780 0.860 7.620 1.100 ;
        RECT  7.490 2.900 7.520 3.140 ;
        RECT  7.250 1.400 7.490 3.140 ;
        RECT  7.090 1.400 7.250 1.640 ;
        RECT  5.020 2.900 7.250 3.140 ;
        RECT  5.890 3.940 6.290 4.250 ;
        RECT  5.540 0.860 5.780 2.620 ;
        RECT  5.300 2.220 5.540 2.620 ;
        RECT  5.020 1.580 5.260 1.820 ;
        RECT  4.780 1.580 5.020 3.140 ;
        RECT  2.220 1.000 4.910 1.240 ;
        RECT  2.510 2.750 4.780 2.990 ;
        RECT  4.150 3.270 4.390 3.660 ;
        RECT  1.890 3.270 4.150 3.510 ;
        RECT  2.270 2.340 2.510 2.990 ;
        RECT  2.150 2.340 2.270 2.580 ;
        RECT  1.980 1.000 2.220 1.570 ;
        RECT  1.910 2.180 2.150 2.580 ;
        RECT  1.630 1.330 1.980 1.570 ;
        RECT  1.650 2.850 1.890 3.750 ;
        RECT  1.630 2.850 1.650 3.090 ;
        RECT  1.390 1.330 1.630 3.090 ;
        RECT  1.110 4.130 1.580 4.370 ;
        RECT  1.110 0.740 1.500 0.980 ;
        RECT  0.870 0.740 1.110 4.370 ;
    END
END TLATSRX2

MACRO TLATSRX1
    CLASS CORE ;
    FOREIGN TLATSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATSRXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.180 1.960 0.190 2.510 ;
        RECT  0.190 1.900 0.200 2.510 ;
        RECT  0.200 1.830 0.460 2.510 ;
        RECT  0.460 1.840 0.510 2.510 ;
        RECT  0.510 1.900 0.590 2.510 ;
        RECT  0.590 1.960 0.600 2.510 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.530 2.090 ;
        RECT  3.530 1.830 3.760 2.620 ;
        RECT  3.760 1.840 3.770 2.620 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  10.650 2.990 10.770 3.390 ;
        RECT  10.760 2.390 10.770 2.650 ;
        RECT  10.650 1.290 10.770 1.830 ;
        RECT  10.770 1.290 11.010 3.390 ;
        RECT  11.010 2.390 11.020 2.650 ;
        RECT  11.010 2.990 11.050 3.390 ;
        RECT  11.010 1.290 11.050 1.950 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.330 2.940 9.570 3.340 ;
        RECT  9.570 2.940 9.580 3.210 ;
        RECT  9.310 1.420 9.580 1.660 ;
        RECT  9.580 1.420 9.700 3.210 ;
        RECT  9.700 1.420 9.820 3.200 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  6.140 1.830 6.150 2.090 ;
        RECT  6.150 1.830 6.400 2.140 ;
        RECT  6.400 1.900 6.520 2.140 ;
        RECT  6.520 1.900 6.920 2.300 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.780 1.950 2.840 2.640 ;
        RECT  2.840 1.950 3.020 2.650 ;
        RECT  3.020 2.390 3.100 2.650 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 3.100 5.440 ;
        RECT  3.100 4.160 3.500 5.440 ;
        RECT  3.500 4.640 6.480 5.440 ;
        RECT  6.480 4.480 6.880 5.440 ;
        RECT  6.880 4.640 8.440 5.440 ;
        RECT  8.440 4.480 8.840 5.440 ;
        RECT  8.840 4.640 10.040 5.440 ;
        RECT  10.040 4.480 10.440 5.440 ;
        RECT  10.440 4.640 11.220 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 2.390 0.400 ;
        RECT  2.390 -0.400 2.790 0.560 ;
        RECT  2.790 -0.400 6.190 0.400 ;
        RECT  6.190 -0.400 6.590 0.560 ;
        RECT  6.590 -0.400 8.480 0.400 ;
        RECT  8.480 -0.400 8.880 1.780 ;
        RECT  8.880 -0.400 10.040 0.400 ;
        RECT  10.040 -0.400 10.440 0.560 ;
        RECT  10.440 -0.400 11.220 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.110 0.880 10.350 4.020 ;
        RECT  9.710 0.880 10.110 1.120 ;
        RECT  9.710 3.780 10.110 4.020 ;
        RECT  9.440 0.670 9.710 1.120 ;
        RECT  9.470 3.780 9.710 4.360 ;
        RECT  9.310 3.940 9.470 4.360 ;
        RECT  9.310 0.670 9.440 0.910 ;
        RECT  6.200 3.940 9.310 4.180 ;
        RECT  8.940 2.060 9.280 2.460 ;
        RECT  8.700 2.060 8.940 3.660 ;
        RECT  4.820 3.420 8.700 3.660 ;
        RECT  7.960 0.680 8.200 3.130 ;
        RECT  7.740 0.680 7.960 1.100 ;
        RECT  7.770 2.890 7.960 3.130 ;
        RECT  5.710 0.860 7.740 1.100 ;
        RECT  7.440 1.870 7.680 2.270 ;
        RECT  7.200 1.390 7.440 3.140 ;
        RECT  6.980 1.390 7.200 1.630 ;
        RECT  4.370 2.900 7.200 3.140 ;
        RECT  5.800 3.940 6.200 4.350 ;
        RECT  5.470 0.860 5.710 2.620 ;
        RECT  4.650 2.380 5.470 2.620 ;
        RECT  4.720 1.580 5.120 1.980 ;
        RECT  4.380 3.420 4.820 3.690 ;
        RECT  2.750 1.010 4.750 1.250 ;
        RECT  4.370 1.740 4.720 1.980 ;
        RECT  1.890 3.450 4.380 3.690 ;
        RECT  4.130 1.740 4.370 3.140 ;
        RECT  3.890 2.900 4.130 3.140 ;
        RECT  3.650 2.900 3.890 3.170 ;
        RECT  2.480 2.930 3.650 3.170 ;
        RECT  2.510 1.010 2.750 1.570 ;
        RECT  1.780 1.330 2.510 1.570 ;
        RECT  2.240 2.670 2.480 3.170 ;
        RECT  2.150 2.670 2.240 2.910 ;
        RECT  1.910 2.330 2.150 2.910 ;
        RECT  1.230 0.690 2.100 0.930 ;
        RECT  1.650 3.190 1.890 3.690 ;
        RECT  1.630 1.330 1.780 2.030 ;
        RECT  1.110 4.070 1.770 4.310 ;
        RECT  1.630 3.190 1.650 3.430 ;
        RECT  1.540 1.330 1.630 3.430 ;
        RECT  1.390 1.790 1.540 3.430 ;
        RECT  1.110 0.690 1.230 1.510 ;
        RECT  0.990 0.690 1.110 4.310 ;
        RECT  0.870 1.270 0.990 4.310 ;
        RECT  0.830 1.270 0.870 1.510 ;
    END
END TLATSRX1

MACRO TLATSXL
    CLASS CORE ;
    FOREIGN TLATSXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.190 1.960 0.200 2.500 ;
        RECT  0.200 1.830 0.460 2.500 ;
        RECT  0.460 2.100 0.590 2.500 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  10.070 1.200 10.100 2.640 ;
        RECT  9.990 2.990 10.110 3.390 ;
        RECT  10.100 1.200 10.110 2.650 ;
        RECT  10.110 1.200 10.310 3.390 ;
        RECT  10.310 2.390 10.350 3.390 ;
        RECT  10.350 2.390 10.360 2.650 ;
        RECT  10.350 2.990 10.390 3.390 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  8.670 2.940 8.910 3.350 ;
        RECT  8.910 2.940 8.920 3.210 ;
        RECT  8.650 1.460 8.920 1.700 ;
        RECT  8.920 1.460 9.040 3.210 ;
        RECT  9.040 1.460 9.160 3.200 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  5.480 1.270 5.490 1.530 ;
        RECT  5.490 1.270 5.740 1.710 ;
        RECT  5.740 1.470 5.810 1.710 ;
        RECT  5.810 1.470 6.050 1.870 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 1.830 2.990 2.090 ;
        RECT  2.990 1.830 3.100 2.270 ;
        RECT  3.100 1.840 3.310 2.270 ;
        RECT  3.310 1.870 3.390 2.270 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 3.180 5.440 ;
        RECT  3.180 4.080 3.420 5.440 ;
        RECT  3.420 4.640 5.920 5.440 ;
        RECT  5.920 4.480 6.320 5.440 ;
        RECT  6.320 4.640 7.780 5.440 ;
        RECT  7.780 4.480 8.180 5.440 ;
        RECT  8.180 4.640 9.380 5.440 ;
        RECT  9.380 4.480 9.780 5.440 ;
        RECT  9.780 4.640 10.560 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 2.460 0.400 ;
        RECT  2.460 -0.400 2.860 0.560 ;
        RECT  2.860 -0.400 5.270 0.400 ;
        RECT  5.270 -0.400 5.670 0.560 ;
        RECT  5.670 -0.400 7.780 0.400 ;
        RECT  7.780 -0.400 8.180 0.560 ;
        RECT  8.180 -0.400 9.380 0.400 ;
        RECT  9.380 -0.400 9.780 0.560 ;
        RECT  9.780 -0.400 10.560 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  9.450 0.880 9.690 4.100 ;
        RECT  9.050 0.880 9.450 1.120 ;
        RECT  8.900 3.860 9.450 4.100 ;
        RECT  8.790 0.680 9.050 1.120 ;
        RECT  8.650 3.860 8.900 4.180 ;
        RECT  8.650 0.680 8.790 0.920 ;
        RECT  5.650 3.940 8.650 4.180 ;
        RECT  8.210 2.040 8.530 2.440 ;
        RECT  8.130 2.040 8.210 3.660 ;
        RECT  7.970 2.150 8.130 3.660 ;
        RECT  1.890 3.420 7.970 3.660 ;
        RECT  7.450 1.020 7.690 3.140 ;
        RECT  6.890 1.020 7.450 1.260 ;
        RECT  4.600 2.900 7.450 3.140 ;
        RECT  6.830 1.630 7.170 2.030 ;
        RECT  6.830 2.380 6.840 2.620 ;
        RECT  6.610 1.630 6.830 2.620 ;
        RECT  6.580 0.870 6.610 2.620 ;
        RECT  6.370 0.870 6.580 1.870 ;
        RECT  5.120 2.380 6.580 2.620 ;
        RECT  6.150 0.870 6.370 1.110 ;
        RECT  5.230 3.940 5.650 4.230 ;
        RECT  4.880 1.550 5.120 2.620 ;
        RECT  3.910 1.550 4.880 1.790 ;
        RECT  4.360 2.200 4.600 3.140 ;
        RECT  4.200 2.200 4.360 2.600 ;
        RECT  2.400 0.950 4.330 1.190 ;
        RECT  3.670 1.550 3.910 3.140 ;
        RECT  2.410 2.900 3.670 3.140 ;
        RECT  2.350 2.490 2.410 3.140 ;
        RECT  2.160 0.950 2.400 1.560 ;
        RECT  2.170 2.030 2.350 3.140 ;
        RECT  2.110 2.030 2.170 2.730 ;
        RECT  1.680 1.320 2.160 1.560 ;
        RECT  1.680 3.080 1.890 3.660 ;
        RECT  1.150 0.760 1.880 1.000 ;
        RECT  1.150 4.070 1.770 4.310 ;
        RECT  1.650 1.320 1.680 3.660 ;
        RECT  1.440 1.320 1.650 3.400 ;
        RECT  0.910 0.760 1.150 4.310 ;
    END
END TLATSXL

MACRO TLATSX4
    CLASS CORE ;
    FOREIGN TLATSX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATSXL ;
    SIZE 14.520 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.270 2.650 ;
        RECT  0.270 1.960 0.460 2.650 ;
        RECT  0.460 1.960 0.510 2.640 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.650 1.820 12.690 3.220 ;
        RECT  12.690 1.230 13.000 3.220 ;
        RECT  13.000 1.230 13.090 3.250 ;
        RECT  13.090 2.850 13.400 3.250 ;
        RECT  13.090 1.230 13.400 1.630 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.330 1.820 11.460 3.220 ;
        RECT  11.460 1.230 11.780 3.250 ;
        RECT  11.780 2.850 11.860 3.250 ;
        RECT  11.780 1.230 11.860 1.630 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  7.420 1.470 7.460 1.870 ;
        RECT  7.460 1.470 7.720 2.090 ;
        RECT  7.720 1.470 7.820 1.870 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 1.830 2.990 2.090 ;
        RECT  2.990 1.830 3.100 2.610 ;
        RECT  3.100 1.840 3.230 2.610 ;
        RECT  3.230 1.950 3.390 2.610 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 3.270 5.440 ;
        RECT  3.270 3.940 3.670 5.440 ;
        RECT  3.670 4.640 7.640 5.440 ;
        RECT  7.640 4.480 8.040 5.440 ;
        RECT  8.040 4.640 9.340 5.440 ;
        RECT  9.340 4.480 9.740 5.440 ;
        RECT  9.740 4.640 10.720 5.440 ;
        RECT  10.720 4.480 11.120 5.440 ;
        RECT  11.120 4.640 12.260 5.440 ;
        RECT  12.260 4.210 12.660 5.440 ;
        RECT  12.660 4.640 13.670 5.440 ;
        RECT  13.670 4.210 14.070 5.440 ;
        RECT  14.070 4.640 14.520 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 2.370 0.400 ;
        RECT  2.370 -0.400 2.770 0.560 ;
        RECT  2.770 -0.400 4.940 0.400 ;
        RECT  4.940 -0.400 5.340 0.560 ;
        RECT  5.340 -0.400 7.030 0.400 ;
        RECT  7.030 -0.400 7.430 0.560 ;
        RECT  7.430 -0.400 9.350 0.400 ;
        RECT  9.350 -0.400 9.750 1.190 ;
        RECT  9.750 -0.400 10.850 0.400 ;
        RECT  10.850 -0.400 11.250 0.950 ;
        RECT  11.250 -0.400 12.260 0.400 ;
        RECT  12.260 -0.400 12.660 0.950 ;
        RECT  12.660 -0.400 13.670 0.400 ;
        RECT  13.670 -0.400 14.070 0.950 ;
        RECT  14.070 -0.400 14.520 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  13.680 2.040 13.920 3.910 ;
        RECT  10.470 3.670 13.680 3.910 ;
        RECT  10.820 1.270 11.060 3.050 ;
        RECT  10.110 1.270 10.820 1.510 ;
        RECT  10.470 2.810 10.820 3.050 ;
        RECT  10.230 2.810 10.470 4.180 ;
        RECT  9.870 2.120 10.300 2.360 ;
        RECT  7.360 3.940 10.230 4.180 ;
        RECT  9.630 2.120 9.870 3.660 ;
        RECT  1.930 3.420 9.630 3.660 ;
        RECT  9.070 2.900 9.130 3.140 ;
        RECT  8.830 0.870 9.070 3.140 ;
        RECT  8.670 0.870 8.830 1.270 ;
        RECT  6.450 2.900 8.830 3.140 ;
        RECT  8.430 1.600 8.550 2.000 ;
        RECT  8.390 1.600 8.430 2.620 ;
        RECT  8.150 0.860 8.390 2.620 ;
        RECT  6.840 0.860 8.150 1.100 ;
        RECT  8.140 1.840 8.150 2.620 ;
        RECT  8.000 2.380 8.140 2.620 ;
        RECT  6.960 3.940 7.360 4.250 ;
        RECT  6.600 0.860 6.840 1.750 ;
        RECT  5.740 1.510 6.600 1.750 ;
        RECT  6.210 2.200 6.450 3.140 ;
        RECT  6.050 2.200 6.210 2.600 ;
        RECT  4.630 0.920 6.090 1.160 ;
        RECT  5.500 1.510 5.740 2.900 ;
        RECT  4.250 2.660 5.500 2.900 ;
        RECT  4.390 0.920 4.630 1.390 ;
        RECT  2.480 1.150 4.390 1.390 ;
        RECT  4.010 2.660 4.250 3.130 ;
        RECT  2.580 2.890 4.010 3.130 ;
        RECT  2.340 2.370 2.580 3.130 ;
        RECT  2.240 1.150 2.480 1.570 ;
        RECT  2.110 2.370 2.340 2.610 ;
        RECT  1.770 1.330 2.240 1.570 ;
        RECT  1.870 2.210 2.110 2.610 ;
        RECT  1.190 0.760 1.960 1.000 ;
        RECT  1.580 2.980 1.930 3.880 ;
        RECT  1.580 1.330 1.770 1.920 ;
        RECT  1.530 1.330 1.580 3.880 ;
        RECT  1.340 1.680 1.530 3.220 ;
        RECT  1.060 0.760 1.190 1.390 ;
        RECT  1.060 3.570 1.170 3.810 ;
        RECT  0.950 0.760 1.060 3.810 ;
        RECT  0.820 1.150 0.950 3.810 ;
        RECT  0.770 1.150 0.820 1.390 ;
        RECT  0.770 3.570 0.820 3.810 ;
    END
END TLATSX4

MACRO TLATSX2
    CLASS CORE ;
    FOREIGN TLATSX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATSXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.310 2.090 ;
        RECT  0.310 1.830 0.460 2.520 ;
        RECT  0.460 1.840 0.550 2.520 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  10.730 0.740 10.970 4.210 ;
        RECT  10.970 2.390 11.010 3.520 ;
        RECT  11.010 2.390 11.020 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  8.780 2.950 9.120 3.210 ;
        RECT  9.120 2.810 9.280 3.210 ;
        RECT  8.950 1.410 9.280 1.650 ;
        RECT  9.280 1.410 9.520 3.210 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  5.480 1.270 5.490 1.530 ;
        RECT  5.490 1.270 5.620 1.710 ;
        RECT  5.620 1.270 5.740 1.990 ;
        RECT  5.740 1.470 5.860 1.990 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 1.830 2.990 2.090 ;
        RECT  2.990 1.830 3.100 2.580 ;
        RECT  3.100 1.840 3.230 2.580 ;
        RECT  3.230 2.180 3.390 2.580 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.790 0.560 5.440 ;
        RECT  0.560 4.640 3.380 5.440 ;
        RECT  3.380 4.080 3.620 5.440 ;
        RECT  3.620 4.640 5.940 5.440 ;
        RECT  5.940 4.480 6.340 5.440 ;
        RECT  6.340 4.640 7.740 5.440 ;
        RECT  7.740 4.480 8.140 5.440 ;
        RECT  8.140 4.640 9.890 5.440 ;
        RECT  9.890 4.190 10.290 5.440 ;
        RECT  10.290 4.640 11.220 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 2.440 0.400 ;
        RECT  2.440 -0.400 2.840 0.560 ;
        RECT  2.840 -0.400 5.190 0.400 ;
        RECT  5.190 -0.400 5.590 0.560 ;
        RECT  5.590 -0.400 7.690 0.400 ;
        RECT  7.690 -0.400 8.090 1.130 ;
        RECT  8.090 -0.400 9.830 0.400 ;
        RECT  9.830 -0.400 10.230 0.560 ;
        RECT  10.230 -0.400 11.220 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.160 0.880 10.400 3.910 ;
        RECT  9.430 0.880 10.160 1.120 ;
        RECT  8.990 3.670 10.160 3.910 ;
        RECT  9.190 0.680 9.430 1.120 ;
        RECT  8.510 0.680 9.190 0.920 ;
        RECT  8.980 3.660 8.990 3.910 ;
        RECT  8.590 3.660 8.980 4.180 ;
        RECT  8.210 2.120 8.700 2.360 ;
        RECT  5.650 3.940 8.590 4.180 ;
        RECT  7.970 2.120 8.210 3.660 ;
        RECT  1.890 3.420 7.970 3.660 ;
        RECT  7.450 1.420 7.690 3.140 ;
        RECT  7.410 1.420 7.450 1.660 ;
        RECT  4.600 2.900 7.450 3.140 ;
        RECT  7.170 0.920 7.410 1.660 ;
        RECT  6.810 0.920 7.170 1.160 ;
        RECT  6.830 1.600 6.890 2.000 ;
        RECT  6.590 1.600 6.830 2.620 ;
        RECT  6.390 1.600 6.590 1.840 ;
        RECT  5.120 2.380 6.590 2.620 ;
        RECT  6.150 0.830 6.390 1.840 ;
        RECT  5.230 3.940 5.650 4.230 ;
        RECT  4.880 1.550 5.120 2.620 ;
        RECT  3.920 1.550 4.880 1.790 ;
        RECT  4.360 2.200 4.600 3.140 ;
        RECT  4.200 2.200 4.360 2.600 ;
        RECT  2.480 0.860 4.250 1.100 ;
        RECT  3.680 1.550 3.920 3.140 ;
        RECT  2.480 2.900 3.680 3.140 ;
        RECT  2.240 0.860 2.480 1.560 ;
        RECT  2.240 2.390 2.480 3.140 ;
        RECT  1.810 1.320 2.240 1.560 ;
        RECT  2.150 2.390 2.240 2.630 ;
        RECT  1.910 2.180 2.150 2.630 ;
        RECT  1.240 0.770 1.960 1.010 ;
        RECT  1.650 2.980 1.890 3.880 ;
        RECT  1.630 1.320 1.810 1.890 ;
        RECT  1.630 2.980 1.650 3.220 ;
        RECT  1.570 1.320 1.630 3.220 ;
        RECT  1.390 1.650 1.570 3.220 ;
        RECT  1.110 0.770 1.240 1.330 ;
        RECT  1.000 0.770 1.110 3.240 ;
        RECT  0.870 1.090 1.000 3.240 ;
        RECT  0.830 1.090 0.870 1.330 ;
    END
END TLATSX2

MACRO TLATSX1
    CLASS CORE ;
    FOREIGN TLATSX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATSXL ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.190 2.040 0.200 2.440 ;
        RECT  0.200 1.830 0.460 2.440 ;
        RECT  0.460 2.010 0.510 2.440 ;
        RECT  0.510 2.040 0.590 2.440 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.990 2.990 10.110 3.390 ;
        RECT  10.100 2.390 10.110 2.650 ;
        RECT  9.990 1.300 10.110 1.830 ;
        RECT  10.110 1.300 10.350 3.390 ;
        RECT  10.350 2.390 10.360 2.650 ;
        RECT  10.350 2.990 10.390 3.390 ;
        RECT  10.350 1.300 10.390 1.960 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  8.590 2.940 8.880 3.340 ;
        RECT  8.650 1.520 8.880 1.760 ;
        RECT  8.880 1.520 8.990 3.340 ;
        RECT  8.990 1.520 9.040 3.210 ;
        RECT  9.040 1.520 9.120 3.200 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  5.390 1.610 6.060 2.100 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.750 1.690 3.270 2.100 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.700 0.560 5.440 ;
        RECT  0.560 4.640 3.100 5.440 ;
        RECT  3.100 4.080 3.500 5.440 ;
        RECT  3.500 4.640 5.930 5.440 ;
        RECT  5.930 4.480 6.330 5.440 ;
        RECT  6.330 4.640 7.780 5.440 ;
        RECT  7.780 4.480 8.180 5.440 ;
        RECT  8.180 4.640 9.380 5.440 ;
        RECT  9.380 4.480 9.780 5.440 ;
        RECT  9.780 4.640 10.560 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 2.500 0.400 ;
        RECT  2.500 -0.400 2.900 0.560 ;
        RECT  2.900 -0.400 5.270 0.400 ;
        RECT  5.270 -0.400 5.670 0.560 ;
        RECT  5.670 -0.400 7.770 0.400 ;
        RECT  7.770 -0.400 8.170 0.560 ;
        RECT  8.170 -0.400 9.380 0.400 ;
        RECT  9.380 -0.400 9.780 0.560 ;
        RECT  9.780 -0.400 10.560 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  9.450 0.880 9.690 4.020 ;
        RECT  9.050 0.880 9.450 1.120 ;
        RECT  9.050 3.780 9.450 4.020 ;
        RECT  8.650 0.670 9.050 1.120 ;
        RECT  8.810 3.780 9.050 4.320 ;
        RECT  8.650 3.940 8.810 4.320 ;
        RECT  5.650 3.940 8.650 4.180 ;
        RECT  8.270 2.040 8.570 2.440 ;
        RECT  8.030 2.040 8.270 3.660 ;
        RECT  1.970 3.420 8.030 3.660 ;
        RECT  7.450 0.870 7.690 3.140 ;
        RECT  7.290 0.870 7.450 1.110 ;
        RECT  4.450 2.900 7.450 3.140 ;
        RECT  6.890 0.690 7.290 1.110 ;
        RECT  6.930 1.460 7.170 2.620 ;
        RECT  6.610 1.460 6.930 1.700 ;
        RECT  5.030 2.380 6.930 2.620 ;
        RECT  6.370 0.910 6.610 1.700 ;
        RECT  6.150 0.910 6.370 1.150 ;
        RECT  5.230 3.940 5.650 4.230 ;
        RECT  4.790 1.630 5.030 2.620 ;
        RECT  4.590 1.630 4.790 1.870 ;
        RECT  4.190 1.470 4.590 1.870 ;
        RECT  4.210 2.200 4.450 3.140 ;
        RECT  3.890 0.780 4.290 1.180 ;
        RECT  3.910 1.630 4.190 1.870 ;
        RECT  3.670 1.630 3.910 2.610 ;
        RECT  2.480 0.940 3.890 1.180 ;
        RECT  2.370 2.370 3.670 2.610 ;
        RECT  2.240 0.940 2.480 1.490 ;
        RECT  2.130 1.990 2.370 2.610 ;
        RECT  1.690 1.250 2.240 1.490 ;
        RECT  1.970 1.990 2.130 2.390 ;
        RECT  1.690 3.020 1.970 3.660 ;
        RECT  1.150 0.700 1.960 0.940 ;
        RECT  1.150 4.010 1.770 4.250 ;
        RECT  1.450 1.250 1.690 3.660 ;
        RECT  0.910 0.700 1.150 4.250 ;
    END
END TLATSX1

MACRO TLATRXL
    CLASS CORE ;
    FOREIGN TLATRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.820 1.640 2.840 2.640 ;
        RECT  2.840 1.640 3.060 2.650 ;
        RECT  3.060 2.370 3.100 2.650 ;
        RECT  3.100 2.370 3.750 2.610 ;
        RECT  3.750 2.370 3.850 2.640 ;
        RECT  3.850 2.370 4.050 2.660 ;
        RECT  4.050 2.370 4.290 2.770 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  8.010 1.180 8.120 1.580 ;
        RECT  8.010 3.040 8.130 3.440 ;
        RECT  8.120 1.180 8.130 2.090 ;
        RECT  8.130 1.180 8.370 3.440 ;
        RECT  8.370 1.180 8.380 2.090 ;
        RECT  8.370 3.040 8.410 3.440 ;
        RECT  8.380 1.180 8.410 1.580 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.570 0.670 6.760 0.910 ;
        RECT  6.750 3.520 6.800 4.010 ;
        RECT  6.800 3.510 6.990 4.010 ;
        RECT  6.760 0.670 7.000 1.100 ;
        RECT  6.990 3.510 7.060 3.770 ;
        RECT  7.060 3.520 7.490 3.760 ;
        RECT  7.000 0.860 7.490 1.100 ;
        RECT  7.490 0.860 7.730 3.760 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.210 2.090 ;
        RECT  0.210 1.830 0.460 2.450 ;
        RECT  0.460 2.050 0.650 2.450 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 2.570 2.190 2.970 ;
        RECT  2.180 1.830 2.190 2.090 ;
        RECT  2.190 1.830 2.430 2.970 ;
        RECT  2.430 1.830 2.440 2.090 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.820 5.440 ;
        RECT  1.820 3.930 2.180 5.440 ;
        RECT  2.180 4.640 3.880 5.440 ;
        RECT  3.880 4.480 4.280 5.440 ;
        RECT  4.280 4.640 5.850 5.440 ;
        RECT  5.850 3.780 6.250 5.440 ;
        RECT  6.250 4.640 7.400 5.440 ;
        RECT  7.400 4.480 7.800 5.440 ;
        RECT  7.800 4.640 8.580 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.970 0.400 ;
        RECT  1.970 -0.400 2.370 0.560 ;
        RECT  2.370 -0.400 5.760 0.400 ;
        RECT  5.760 -0.400 6.000 1.140 ;
        RECT  6.000 -0.400 7.310 0.400 ;
        RECT  7.310 -0.400 7.710 0.560 ;
        RECT  7.710 -0.400 8.580 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.970 1.460 7.210 3.180 ;
        RECT  6.580 1.460 6.970 1.700 ;
        RECT  6.670 2.720 6.970 3.180 ;
        RECT  5.770 2.720 6.670 2.960 ;
        RECT  6.170 2.040 6.570 2.440 ;
        RECT  5.250 2.120 6.170 2.360 ;
        RECT  5.530 2.640 5.770 3.040 ;
        RECT  5.010 0.700 5.250 4.120 ;
        RECT  3.880 0.700 5.010 0.940 ;
        RECT  3.540 3.880 5.010 4.120 ;
        RECT  4.490 3.100 4.730 3.500 ;
        RECT  1.820 3.260 4.490 3.500 ;
        RECT  3.580 1.270 3.860 1.510 ;
        RECT  3.340 0.870 3.580 1.510 ;
        RECT  3.140 3.780 3.540 4.180 ;
        RECT  1.820 0.870 3.340 1.110 ;
        RECT  1.580 0.870 1.820 3.660 ;
        RECT  1.480 0.870 1.580 1.110 ;
        RECT  1.320 3.410 1.580 3.660 ;
        RECT  1.160 0.730 1.480 1.110 ;
        RECT  1.000 3.410 1.320 3.940 ;
        RECT  1.230 2.240 1.290 2.640 ;
        RECT  1.150 1.460 1.230 3.140 ;
        RECT  1.080 0.730 1.160 0.970 ;
        RECT  0.990 1.380 1.150 3.140 ;
        RECT  0.920 3.540 1.000 3.940 ;
        RECT  0.910 1.380 0.990 1.780 ;
        RECT  0.830 2.900 0.990 3.140 ;
    END
END TLATRXL

MACRO TLATRX4
    CLASS CORE ;
    FOREIGN TLATRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATRXL ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.770 2.380 3.200 2.930 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  10.670 1.260 10.700 2.660 ;
        RECT  10.700 1.220 10.710 2.660 ;
        RECT  10.710 1.220 11.100 3.210 ;
        RECT  11.100 1.260 11.110 3.210 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.120 1.760 9.300 3.210 ;
        RECT  9.300 1.420 9.310 3.210 ;
        RECT  9.310 1.220 9.520 3.210 ;
        RECT  9.520 1.220 9.710 2.660 ;
        RECT  9.710 1.260 9.790 2.660 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  5.480 1.710 6.130 2.110 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.720 2.090 ;
        RECT  1.720 1.830 1.780 2.460 ;
        RECT  1.780 1.840 1.960 2.460 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 2.730 5.440 ;
        RECT  2.730 4.480 3.130 5.440 ;
        RECT  3.130 4.640 4.950 5.440 ;
        RECT  4.950 4.480 5.350 5.440 ;
        RECT  5.350 4.640 7.100 5.440 ;
        RECT  7.100 4.480 7.500 5.440 ;
        RECT  7.500 4.640 8.320 5.440 ;
        RECT  8.320 4.480 8.720 5.440 ;
        RECT  8.720 4.640 9.860 5.440 ;
        RECT  9.860 4.090 10.260 5.440 ;
        RECT  10.260 4.640 11.440 5.440 ;
        RECT  11.440 4.090 11.840 5.440 ;
        RECT  11.840 4.640 12.540 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 2.030 0.400 ;
        RECT  2.030 -0.400 2.430 1.010 ;
        RECT  2.430 -0.400 5.570 0.400 ;
        RECT  5.570 -0.400 5.970 0.560 ;
        RECT  5.970 -0.400 8.510 0.400 ;
        RECT  8.510 -0.400 8.910 0.560 ;
        RECT  8.910 -0.400 10.050 0.400 ;
        RECT  10.050 -0.400 10.450 0.940 ;
        RECT  10.450 -0.400 11.310 0.400 ;
        RECT  11.310 -0.400 11.710 0.940 ;
        RECT  11.710 -0.400 12.540 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  11.380 1.790 11.620 3.730 ;
        RECT  8.870 3.490 11.380 3.730 ;
        RECT  8.630 1.620 8.870 3.730 ;
        RECT  8.390 1.620 8.630 1.860 ;
        RECT  8.210 3.490 8.630 3.730 ;
        RECT  7.990 1.460 8.390 1.860 ;
        RECT  8.110 2.170 8.350 2.780 ;
        RECT  7.970 3.080 8.210 4.180 ;
        RECT  7.730 2.540 8.110 2.780 ;
        RECT  4.670 3.940 7.970 4.180 ;
        RECT  7.490 2.540 7.730 3.660 ;
        RECT  7.280 1.230 7.650 1.630 ;
        RECT  1.850 3.420 7.490 3.660 ;
        RECT  7.240 0.860 7.280 1.630 ;
        RECT  7.040 0.860 7.240 3.140 ;
        RECT  5.120 0.860 7.040 1.100 ;
        RECT  7.000 1.390 7.040 3.140 ;
        RECT  6.320 2.900 7.000 3.140 ;
        RECT  6.520 1.380 6.760 2.620 ;
        RECT  6.430 1.380 6.520 1.780 ;
        RECT  6.050 2.380 6.520 2.620 ;
        RECT  5.810 2.380 6.050 3.140 ;
        RECT  3.710 2.900 5.810 3.140 ;
        RECT  4.880 0.860 5.120 2.560 ;
        RECT  3.990 2.320 4.880 2.560 ;
        RECT  4.270 3.940 4.670 4.230 ;
        RECT  3.710 1.600 4.500 1.840 ;
        RECT  3.050 1.030 4.170 1.270 ;
        RECT  3.550 3.940 3.950 4.230 ;
        RECT  3.470 1.600 3.710 3.140 ;
        RECT  2.430 3.940 3.550 4.180 ;
        RECT  3.450 1.600 3.470 2.110 ;
        RECT  2.480 1.870 3.450 2.110 ;
        RECT  2.810 1.030 3.050 1.580 ;
        RECT  1.060 1.290 2.810 1.580 ;
        RECT  2.240 1.870 2.480 3.100 ;
        RECT  2.190 3.940 2.430 4.370 ;
        RECT  1.380 2.860 2.240 3.100 ;
        RECT  1.130 4.130 2.190 4.370 ;
        RECT  1.450 3.420 1.850 3.850 ;
        RECT  1.060 3.420 1.450 3.660 ;
        RECT  0.890 3.940 1.130 4.370 ;
        RECT  0.820 1.290 1.060 3.660 ;
        RECT  0.500 3.940 0.890 4.180 ;
        RECT  0.570 1.290 0.820 1.670 ;
        RECT  0.170 0.770 0.570 1.670 ;
        RECT  0.260 1.910 0.500 4.180 ;
    END
END TLATRX4

MACRO TLATRX2
    CLASS CORE ;
    FOREIGN TLATRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATRXL ;
    SIZE 9.240 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.040 2.310 3.200 2.710 ;
        RECT  3.200 2.310 3.440 3.130 ;
        RECT  3.440 2.890 4.160 3.130 ;
        RECT  4.160 2.890 4.420 3.210 ;
        RECT  4.420 2.890 4.520 3.200 ;
        RECT  4.520 2.890 4.600 3.130 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  8.120 3.510 8.140 3.770 ;
        RECT  8.140 3.500 8.380 3.770 ;
        RECT  8.380 3.500 8.650 3.740 ;
        RECT  8.650 1.380 8.790 1.780 ;
        RECT  8.650 2.910 8.830 3.740 ;
        RECT  8.790 1.380 8.830 1.840 ;
        RECT  8.830 1.380 8.890 3.740 ;
        RECT  8.890 1.380 9.070 3.520 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  7.300 2.960 7.350 4.250 ;
        RECT  7.350 1.390 7.540 4.250 ;
        RECT  7.540 1.390 7.590 3.210 ;
        RECT  7.590 2.950 7.720 3.210 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.460 2.450 ;
        RECT  0.460 2.050 0.600 2.450 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 2.390 2.190 2.650 ;
        RECT  2.190 2.390 2.260 2.710 ;
        RECT  2.260 2.300 2.580 2.710 ;
        RECT  2.580 2.300 2.660 2.700 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.790 5.440 ;
        RECT  1.790 4.230 2.190 5.440 ;
        RECT  2.190 4.640 3.880 5.440 ;
        RECT  3.880 4.480 4.280 5.440 ;
        RECT  4.280 4.640 5.970 5.440 ;
        RECT  5.970 4.480 6.370 5.440 ;
        RECT  6.370 4.640 8.040 5.440 ;
        RECT  8.040 4.110 8.440 5.440 ;
        RECT  8.440 4.640 9.240 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 2.210 0.400 ;
        RECT  2.210 -0.400 2.610 0.560 ;
        RECT  2.610 -0.400 5.750 0.400 ;
        RECT  5.750 -0.400 6.150 0.560 ;
        RECT  6.150 -0.400 7.980 0.400 ;
        RECT  7.980 -0.400 8.380 0.560 ;
        RECT  8.380 -0.400 9.240 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  8.320 2.070 8.550 2.470 ;
        RECT  8.310 0.860 8.320 2.470 ;
        RECT  8.080 0.860 8.310 2.310 ;
        RECT  7.020 0.860 8.080 1.100 ;
        RECT  6.860 0.680 7.020 3.310 ;
        RECT  6.780 0.680 6.860 3.390 ;
        RECT  6.620 0.680 6.780 1.990 ;
        RECT  6.620 2.990 6.780 3.390 ;
        RECT  6.610 0.680 6.620 1.100 ;
        RECT  6.160 1.590 6.620 1.990 ;
        RECT  5.860 2.310 6.490 2.710 ;
        RECT  5.620 0.860 5.860 4.180 ;
        RECT  5.250 0.860 5.620 1.100 ;
        RECT  3.410 3.940 5.620 4.180 ;
        RECT  5.150 3.340 5.320 3.580 ;
        RECT  5.010 0.680 5.250 1.100 ;
        RECT  4.910 2.240 5.150 3.580 ;
        RECT  4.030 0.680 5.010 0.920 ;
        RECT  4.160 2.240 4.910 2.480 ;
        RECT  4.700 1.680 4.880 1.920 ;
        RECT  4.460 1.200 4.700 1.920 ;
        RECT  2.530 1.200 4.460 1.440 ;
        RECT  3.920 1.730 4.160 2.480 ;
        RECT  1.980 1.730 3.920 1.970 ;
        RECT  3.010 3.860 3.410 4.180 ;
        RECT  2.290 0.860 2.530 1.440 ;
        RECT  1.160 0.860 2.290 1.100 ;
        RECT  1.820 1.380 1.980 1.970 ;
        RECT  1.580 1.380 1.820 3.900 ;
        RECT  1.310 3.660 1.580 3.900 ;
        RECT  0.910 3.660 1.310 4.060 ;
        RECT  1.160 2.030 1.300 2.430 ;
        RECT  1.120 0.860 1.160 2.430 ;
        RECT  0.920 0.860 1.120 3.150 ;
        RECT  0.880 2.170 0.920 3.150 ;
    END
END TLATRX2

MACRO TLATRX1
    CLASS CORE ;
    FOREIGN TLATRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATRXL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.410 2.900 3.570 3.140 ;
        RECT  3.570 2.410 3.810 3.140 ;
        RECT  3.810 2.410 4.160 2.650 ;
        RECT  4.160 2.390 4.320 2.650 ;
        RECT  4.320 2.090 4.560 2.650 ;
        RECT  4.560 2.090 5.150 2.330 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  8.010 1.170 8.120 1.830 ;
        RECT  8.010 2.930 8.130 3.330 ;
        RECT  8.120 1.170 8.130 2.090 ;
        RECT  8.130 1.170 8.370 3.330 ;
        RECT  8.370 1.170 8.380 2.090 ;
        RECT  8.370 2.930 8.410 3.330 ;
        RECT  8.380 1.170 8.410 1.960 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.550 0.670 6.790 0.910 ;
        RECT  6.750 3.520 6.800 4.170 ;
        RECT  6.800 3.510 6.990 4.170 ;
        RECT  6.790 0.670 7.030 1.100 ;
        RECT  6.990 3.510 7.060 3.770 ;
        RECT  7.060 3.520 7.490 3.760 ;
        RECT  7.030 0.860 7.490 1.100 ;
        RECT  7.490 0.860 7.730 3.760 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.180 2.070 0.200 2.470 ;
        RECT  0.200 1.830 0.460 2.470 ;
        RECT  0.460 2.070 0.580 2.470 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.110 2.400 2.180 3.120 ;
        RECT  2.180 2.390 2.280 3.120 ;
        RECT  2.280 1.700 2.520 3.120 ;
        RECT  2.520 1.700 2.770 1.940 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.930 5.440 ;
        RECT  1.930 3.940 2.170 5.440 ;
        RECT  2.170 4.640 3.970 5.440 ;
        RECT  3.970 4.480 4.370 5.440 ;
        RECT  4.370 4.640 5.870 5.440 ;
        RECT  5.870 4.070 6.270 5.440 ;
        RECT  6.270 4.640 7.400 5.440 ;
        RECT  7.400 4.480 7.800 5.440 ;
        RECT  7.800 4.640 8.580 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 2.100 0.400 ;
        RECT  2.100 -0.400 2.500 0.560 ;
        RECT  2.500 -0.400 5.890 0.400 ;
        RECT  5.890 -0.400 6.130 0.880 ;
        RECT  6.130 -0.400 7.310 0.400 ;
        RECT  7.310 -0.400 7.710 0.560 ;
        RECT  7.710 -0.400 8.580 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.970 1.460 7.210 3.180 ;
        RECT  6.630 1.460 6.970 1.700 ;
        RECT  6.670 2.780 6.970 3.180 ;
        RECT  6.400 2.940 6.670 3.180 ;
        RECT  6.170 2.040 6.570 2.440 ;
        RECT  6.160 2.940 6.400 3.370 ;
        RECT  5.630 2.120 6.170 2.360 ;
        RECT  5.500 3.130 6.160 3.370 ;
        RECT  5.390 1.000 5.630 2.850 ;
        RECT  3.910 1.000 5.390 1.240 ;
        RECT  5.220 2.610 5.390 2.850 ;
        RECT  4.980 2.610 5.220 3.880 ;
        RECT  4.890 3.640 4.980 3.880 ;
        RECT  4.610 3.640 4.890 4.180 ;
        RECT  4.330 2.940 4.700 3.340 ;
        RECT  3.470 3.940 4.610 4.180 ;
        RECT  4.300 2.940 4.330 3.660 ;
        RECT  4.090 3.080 4.300 3.660 ;
        RECT  3.100 3.420 4.090 3.660 ;
        RECT  3.290 1.740 3.990 1.980 ;
        RECT  3.070 3.940 3.470 4.340 ;
        RECT  3.100 1.740 3.290 2.460 ;
        RECT  3.050 1.740 3.100 3.660 ;
        RECT  2.860 2.220 3.050 3.660 ;
        RECT  1.820 3.420 2.860 3.660 ;
        RECT  1.760 1.720 1.820 3.660 ;
        RECT  1.640 0.730 1.760 3.660 ;
        RECT  1.580 0.730 1.640 4.020 ;
        RECT  1.520 0.730 1.580 1.960 ;
        RECT  1.420 3.420 1.580 4.020 ;
        RECT  1.360 0.730 1.520 0.970 ;
        RECT  1.400 3.420 1.420 4.100 ;
        RECT  1.020 3.700 1.400 4.100 ;
        RECT  1.150 2.240 1.300 2.640 ;
        RECT  1.100 1.380 1.150 2.640 ;
        RECT  0.910 1.380 1.100 3.210 ;
        RECT  0.860 2.320 0.910 3.210 ;
    END
END TLATRX1

MACRO TLATNSRXL
    CLASS CORE ;
    FOREIGN TLATNSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.190 2.060 0.200 2.460 ;
        RECT  0.200 1.830 0.460 2.460 ;
        RECT  0.460 2.060 0.590 2.460 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.540 2.090 ;
        RECT  3.540 1.830 3.760 2.590 ;
        RECT  3.760 1.840 3.780 2.590 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  10.650 2.990 10.770 3.390 ;
        RECT  10.760 2.390 10.770 2.650 ;
        RECT  10.650 1.240 10.770 1.830 ;
        RECT  10.770 1.240 11.010 3.390 ;
        RECT  11.010 2.390 11.020 2.650 ;
        RECT  11.010 2.990 11.050 3.390 ;
        RECT  11.010 1.240 11.050 1.960 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.330 2.940 9.570 3.350 ;
        RECT  9.570 2.940 9.580 3.210 ;
        RECT  9.250 1.440 9.580 1.680 ;
        RECT  9.580 1.440 9.700 3.210 ;
        RECT  9.700 1.440 9.820 3.200 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  6.140 1.830 6.150 2.090 ;
        RECT  6.150 1.830 6.400 2.140 ;
        RECT  6.400 1.900 6.520 2.140 ;
        RECT  6.520 1.900 6.920 2.300 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.730 1.940 2.750 2.180 ;
        RECT  2.750 1.940 2.840 2.620 ;
        RECT  2.840 1.940 3.100 2.650 ;
        RECT  3.100 1.940 3.130 2.520 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 3.100 5.440 ;
        RECT  3.100 4.080 3.500 5.440 ;
        RECT  3.500 4.640 6.510 5.440 ;
        RECT  6.510 4.480 6.910 5.440 ;
        RECT  6.910 4.640 8.430 5.440 ;
        RECT  8.430 4.480 8.830 5.440 ;
        RECT  8.830 4.640 10.040 5.440 ;
        RECT  10.040 4.480 10.440 5.440 ;
        RECT  10.440 4.640 11.220 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 2.580 0.400 ;
        RECT  2.580 -0.400 2.980 0.560 ;
        RECT  2.980 -0.400 6.130 0.400 ;
        RECT  6.130 -0.400 6.530 0.560 ;
        RECT  6.530 -0.400 8.360 0.400 ;
        RECT  8.360 -0.400 8.370 1.660 ;
        RECT  8.370 -0.400 8.770 1.780 ;
        RECT  8.770 -0.400 8.780 1.660 ;
        RECT  8.780 -0.400 9.980 0.400 ;
        RECT  9.980 -0.400 10.380 0.560 ;
        RECT  10.380 -0.400 11.220 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.110 0.880 10.350 4.020 ;
        RECT  9.650 0.880 10.110 1.120 ;
        RECT  9.710 3.780 10.110 4.020 ;
        RECT  9.470 3.780 9.710 4.360 ;
        RECT  9.380 0.680 9.650 1.120 ;
        RECT  9.310 3.940 9.470 4.360 ;
        RECT  9.250 0.680 9.380 0.920 ;
        RECT  6.230 3.940 9.310 4.180 ;
        RECT  8.950 2.060 9.230 2.460 ;
        RECT  8.710 2.060 8.950 3.660 ;
        RECT  4.730 3.420 8.710 3.660 ;
        RECT  8.090 2.900 8.170 3.140 ;
        RECT  7.850 0.680 8.090 3.140 ;
        RECT  7.660 0.680 7.850 1.100 ;
        RECT  7.770 2.900 7.850 3.140 ;
        RECT  5.620 0.860 7.660 1.100 ;
        RECT  7.460 1.870 7.570 2.270 ;
        RECT  7.220 1.370 7.460 3.070 ;
        RECT  7.180 1.370 7.220 1.620 ;
        RECT  5.530 2.830 7.220 3.070 ;
        RECT  7.000 1.370 7.180 1.610 ;
        RECT  5.830 3.940 6.230 4.350 ;
        RECT  5.380 0.860 5.620 1.840 ;
        RECT  5.290 2.480 5.530 3.070 ;
        RECT  5.070 1.600 5.380 1.840 ;
        RECT  5.110 2.480 5.290 2.720 ;
        RECT  4.710 2.320 5.110 2.720 ;
        RECT  4.670 1.600 5.070 2.000 ;
        RECT  2.960 1.080 4.810 1.320 ;
        RECT  4.410 3.420 4.730 3.690 ;
        RECT  4.420 1.760 4.670 2.000 ;
        RECT  4.180 1.760 4.420 3.140 ;
        RECT  1.890 3.450 4.410 3.690 ;
        RECT  4.070 2.900 4.180 3.140 ;
        RECT  3.830 2.900 4.070 3.170 ;
        RECT  2.480 2.930 3.830 3.170 ;
        RECT  2.720 1.080 2.960 1.540 ;
        RECT  1.810 1.300 2.720 1.540 ;
        RECT  2.240 2.460 2.480 3.170 ;
        RECT  1.230 0.730 2.290 0.970 ;
        RECT  2.150 2.460 2.240 2.700 ;
        RECT  1.910 2.280 2.150 2.700 ;
        RECT  1.650 2.980 1.890 3.690 ;
        RECT  1.630 1.300 1.810 1.960 ;
        RECT  1.230 4.070 1.770 4.310 ;
        RECT  1.630 2.980 1.650 3.220 ;
        RECT  1.570 1.300 1.630 3.220 ;
        RECT  1.390 1.720 1.570 3.220 ;
        RECT  1.110 0.730 1.230 1.450 ;
        RECT  1.110 3.550 1.230 4.310 ;
        RECT  0.990 0.730 1.110 4.310 ;
        RECT  0.870 1.210 0.990 3.790 ;
        RECT  0.830 1.210 0.870 1.450 ;
        RECT  0.830 3.550 0.870 3.790 ;
    END
END TLATNSRXL

MACRO TLATNSRX4
    CLASS CORE ;
    FOREIGN TLATNSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNSRXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.530 1.780 1.140 2.180 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.780 1.830 8.810 2.090 ;
        RECT  8.810 1.830 9.040 2.310 ;
        RECT  9.040 1.840 9.130 2.310 ;
        RECT  9.130 1.910 9.210 2.310 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.290 1.820 15.390 3.220 ;
        RECT  15.390 1.310 15.500 3.220 ;
        RECT  15.500 1.230 15.640 3.220 ;
        RECT  15.640 1.230 15.730 3.250 ;
        RECT  15.730 2.850 16.040 3.250 ;
        RECT  15.730 1.230 16.040 1.830 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.970 1.820 14.100 3.220 ;
        RECT  14.100 1.230 14.420 3.250 ;
        RECT  14.420 2.850 14.500 3.250 ;
        RECT  14.420 1.230 14.500 1.630 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  10.010 1.480 10.090 1.880 ;
        RECT  10.090 1.480 10.100 2.080 ;
        RECT  10.100 1.480 10.360 2.090 ;
        RECT  10.360 1.480 10.410 1.880 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.510 2.090 ;
        RECT  3.510 1.830 3.750 2.620 ;
        RECT  3.750 1.830 3.760 2.090 ;
        RECT  3.750 2.380 5.270 2.620 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.930 5.440 ;
        RECT  0.930 3.220 1.330 5.440 ;
        RECT  1.330 4.640 6.350 5.440 ;
        RECT  6.350 4.480 6.750 5.440 ;
        RECT  6.750 4.640 9.990 5.440 ;
        RECT  9.990 4.480 10.390 5.440 ;
        RECT  10.390 4.640 11.900 5.440 ;
        RECT  11.900 4.480 12.300 5.440 ;
        RECT  12.300 4.640 13.360 5.440 ;
        RECT  13.360 4.480 13.760 5.440 ;
        RECT  13.760 4.640 14.770 5.440 ;
        RECT  14.770 4.210 15.170 5.440 ;
        RECT  15.170 4.640 16.310 5.440 ;
        RECT  16.310 4.210 16.710 5.440 ;
        RECT  16.710 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.200 0.400 ;
        RECT  1.200 -0.400 1.600 0.560 ;
        RECT  1.600 -0.400 2.960 0.400 ;
        RECT  2.960 -0.400 3.360 0.560 ;
        RECT  3.360 -0.400 5.870 0.400 ;
        RECT  5.870 -0.400 6.270 0.870 ;
        RECT  6.270 -0.400 9.570 0.400 ;
        RECT  9.570 -0.400 9.970 0.560 ;
        RECT  9.970 -0.400 11.990 0.400 ;
        RECT  11.990 -0.400 12.390 0.560 ;
        RECT  12.390 -0.400 13.440 0.400 ;
        RECT  13.440 -0.400 13.840 0.560 ;
        RECT  13.840 -0.400 14.770 0.400 ;
        RECT  14.770 -0.400 15.170 0.950 ;
        RECT  15.170 -0.400 16.310 0.400 ;
        RECT  16.310 -0.400 16.710 0.950 ;
        RECT  16.710 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.400 2.040 16.640 3.860 ;
        RECT  13.030 3.620 16.400 3.860 ;
        RECT  13.460 1.390 13.700 3.020 ;
        RECT  13.000 1.390 13.460 1.630 ;
        RECT  13.030 2.780 13.460 3.020 ;
        RECT  12.450 2.130 13.180 2.370 ;
        RECT  12.790 2.770 13.030 4.180 ;
        RECT  12.600 1.230 13.000 1.630 ;
        RECT  9.710 3.940 12.790 4.180 ;
        RECT  12.210 2.130 12.450 3.660 ;
        RECT  2.550 3.420 12.210 3.660 ;
        RECT  11.680 1.160 11.920 3.140 ;
        RECT  11.500 1.160 11.680 1.400 ;
        RECT  8.410 2.900 11.680 3.140 ;
        RECT  11.260 0.940 11.500 1.400 ;
        RECT  10.980 1.680 11.360 2.080 ;
        RECT  10.960 0.860 10.980 2.080 ;
        RECT  10.740 0.860 10.960 2.620 ;
        RECT  8.800 0.860 10.740 1.100 ;
        RECT  10.720 1.840 10.740 2.620 ;
        RECT  10.550 2.380 10.720 2.620 ;
        RECT  9.390 3.940 9.710 4.230 ;
        RECT  9.310 3.990 9.390 4.230 ;
        RECT  7.430 4.130 8.990 4.370 ;
        RECT  8.560 0.860 8.800 1.480 ;
        RECT  7.770 1.240 8.560 1.480 ;
        RECT  8.170 1.760 8.410 3.140 ;
        RECT  3.080 2.900 8.170 3.140 ;
        RECT  6.950 0.720 8.070 0.960 ;
        RECT  7.530 1.240 7.770 2.600 ;
        RECT  7.370 1.830 7.530 2.600 ;
        RECT  7.190 3.940 7.430 4.370 ;
        RECT  7.350 1.830 7.370 2.520 ;
        RECT  4.150 1.830 7.350 2.070 ;
        RECT  5.990 3.940 7.190 4.180 ;
        RECT  6.710 0.720 6.950 1.390 ;
        RECT  5.530 1.150 6.710 1.390 ;
        RECT  5.750 3.940 5.990 4.360 ;
        RECT  1.870 4.120 5.750 4.360 ;
        RECT  5.290 1.040 5.530 1.390 ;
        RECT  2.550 1.040 5.290 1.280 ;
        RECT  2.840 2.180 3.080 3.140 ;
        RECT  2.310 1.040 2.550 3.660 ;
        RECT  2.150 1.040 2.310 1.450 ;
        RECT  1.870 1.780 2.030 2.180 ;
        RECT  1.630 1.200 1.870 4.360 ;
        RECT  0.630 1.200 1.630 1.440 ;
        RECT  0.570 2.740 1.630 2.980 ;
        RECT  0.230 0.640 0.630 1.540 ;
        RECT  0.250 2.740 0.570 4.300 ;
        RECT  0.170 2.900 0.250 4.300 ;
    END
END TLATNSRX4

MACRO TLATNSRX2
    CLASS CORE ;
    FOREIGN TLATNSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNSRXL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.460 3.020 ;
        RECT  0.460 2.400 0.540 3.020 ;
        RECT  0.540 2.550 0.550 3.020 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.700 1.960 3.860 2.360 ;
        RECT  3.860 1.850 4.100 2.360 ;
        RECT  4.100 1.850 4.160 2.090 ;
        RECT  4.160 1.830 4.420 2.090 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.380 1.370 11.390 3.020 ;
        RECT  11.390 1.200 11.670 3.390 ;
        RECT  11.670 2.390 11.680 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.440 2.950 9.700 3.210 ;
        RECT  9.720 1.410 10.010 1.650 ;
        RECT  9.700 2.960 10.050 3.200 ;
        RECT  10.010 1.410 10.050 1.820 ;
        RECT  10.050 1.410 10.290 3.310 ;
        RECT  10.290 2.910 10.450 3.310 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  6.140 1.830 6.400 2.090 ;
        RECT  6.400 1.850 6.420 2.090 ;
        RECT  6.420 1.850 6.660 2.610 ;
        RECT  6.660 2.370 6.950 2.610 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 1.830 2.980 2.090 ;
        RECT  2.980 1.830 3.100 2.360 ;
        RECT  3.100 1.840 3.380 2.360 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 3.250 5.440 ;
        RECT  3.250 3.790 3.650 5.440 ;
        RECT  3.650 4.640 6.560 5.440 ;
        RECT  6.560 4.480 6.960 5.440 ;
        RECT  6.960 4.640 8.470 5.440 ;
        RECT  8.470 4.480 8.870 5.440 ;
        RECT  8.870 4.640 10.700 5.440 ;
        RECT  10.700 4.190 11.100 5.440 ;
        RECT  11.100 4.640 11.880 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.870 ;
        RECT  0.570 -0.400 2.500 0.400 ;
        RECT  2.500 -0.400 2.900 0.560 ;
        RECT  2.900 -0.400 6.460 0.400 ;
        RECT  6.460 -0.400 6.860 0.560 ;
        RECT  6.860 -0.400 8.450 0.400 ;
        RECT  8.450 -0.400 8.850 0.560 ;
        RECT  8.850 -0.400 10.600 0.400 ;
        RECT  10.600 -0.400 11.000 0.560 ;
        RECT  11.000 -0.400 11.880 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.820 0.880 11.060 3.910 ;
        RECT  9.750 0.880 10.820 1.120 ;
        RECT  9.880 3.670 10.820 3.910 ;
        RECT  9.640 3.670 9.880 4.180 ;
        RECT  9.510 0.670 9.750 1.120 ;
        RECT  6.290 3.940 9.640 4.180 ;
        RECT  9.180 0.670 9.510 0.910 ;
        RECT  9.080 2.040 9.290 2.440 ;
        RECT  8.840 2.040 9.080 3.660 ;
        RECT  4.390 3.420 8.840 3.660 ;
        RECT  8.310 0.860 8.550 3.140 ;
        RECT  8.060 0.860 8.310 1.100 ;
        RECT  7.860 2.900 8.310 3.140 ;
        RECT  7.660 0.670 8.060 1.100 ;
        RECT  7.570 1.900 8.030 2.300 ;
        RECT  5.760 0.860 7.660 1.100 ;
        RECT  7.330 1.410 7.570 3.140 ;
        RECT  7.130 1.410 7.330 1.650 ;
        RECT  5.540 2.900 7.330 3.140 ;
        RECT  5.890 3.940 6.290 4.250 ;
        RECT  5.520 0.860 5.760 1.820 ;
        RECT  5.300 2.220 5.540 3.140 ;
        RECT  5.020 1.580 5.520 1.820 ;
        RECT  4.430 1.000 5.060 1.240 ;
        RECT  4.780 1.580 5.020 2.990 ;
        RECT  2.480 2.750 4.780 2.990 ;
        RECT  4.190 1.000 4.430 1.500 ;
        RECT  4.150 3.270 4.390 3.660 ;
        RECT  2.070 1.260 4.190 1.500 ;
        RECT  1.950 3.270 4.150 3.510 ;
        RECT  2.240 2.340 2.480 2.990 ;
        RECT  2.140 2.340 2.240 2.580 ;
        RECT  1.900 2.180 2.140 2.580 ;
        RECT  1.670 1.180 2.070 1.590 ;
        RECT  1.610 2.860 1.950 3.760 ;
        RECT  1.610 1.350 1.670 1.590 ;
        RECT  1.550 1.350 1.610 3.760 ;
        RECT  1.370 1.350 1.550 3.120 ;
        RECT  1.090 0.670 1.330 1.070 ;
        RECT  0.850 0.670 1.090 3.950 ;
    END
END TLATNSRX2

MACRO TLATNSRX1
    CLASS CORE ;
    FOREIGN TLATNSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNSRXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.260 0.550 2.660 ;
        RECT  0.550 2.090 0.630 2.490 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.530 2.090 ;
        RECT  3.530 1.830 3.760 2.570 ;
        RECT  3.760 1.840 3.770 2.570 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  10.650 1.290 10.670 1.690 ;
        RECT  10.650 2.990 10.770 3.390 ;
        RECT  10.760 2.390 10.770 2.650 ;
        RECT  10.670 1.290 10.770 1.820 ;
        RECT  10.770 1.290 11.010 3.390 ;
        RECT  11.010 2.390 11.020 2.650 ;
        RECT  11.010 2.990 11.050 3.390 ;
        RECT  11.010 1.290 11.050 1.950 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.330 2.940 9.570 3.340 ;
        RECT  9.570 2.940 9.580 3.210 ;
        RECT  9.310 1.420 9.580 1.660 ;
        RECT  9.580 1.420 9.700 3.210 ;
        RECT  9.700 1.420 9.820 3.200 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  6.140 1.830 6.150 2.090 ;
        RECT  6.150 1.830 6.400 2.140 ;
        RECT  6.400 1.900 6.520 2.140 ;
        RECT  6.520 1.900 6.920 2.300 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.800 1.890 2.840 2.640 ;
        RECT  2.840 1.890 3.040 2.650 ;
        RECT  3.040 2.390 3.100 2.650 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 3.100 5.440 ;
        RECT  3.100 4.160 3.500 5.440 ;
        RECT  3.500 4.640 6.480 5.440 ;
        RECT  6.480 4.480 6.880 5.440 ;
        RECT  6.880 4.640 8.440 5.440 ;
        RECT  8.440 4.480 8.840 5.440 ;
        RECT  8.840 4.640 10.040 5.440 ;
        RECT  10.040 4.480 10.440 5.440 ;
        RECT  10.440 4.640 11.220 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 2.470 0.400 ;
        RECT  2.470 -0.400 2.870 0.560 ;
        RECT  2.870 -0.400 6.140 0.400 ;
        RECT  6.140 -0.400 6.540 0.560 ;
        RECT  6.540 -0.400 8.480 0.400 ;
        RECT  8.480 -0.400 8.880 1.790 ;
        RECT  8.880 -0.400 10.040 0.400 ;
        RECT  10.040 -0.400 10.440 0.560 ;
        RECT  10.440 -0.400 11.220 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.110 0.880 10.350 4.020 ;
        RECT  9.710 0.880 10.110 1.120 ;
        RECT  9.710 3.780 10.110 4.020 ;
        RECT  9.450 0.680 9.710 1.120 ;
        RECT  9.470 3.780 9.710 4.370 ;
        RECT  9.310 3.940 9.470 4.370 ;
        RECT  9.310 0.680 9.450 0.920 ;
        RECT  6.200 3.940 9.310 4.180 ;
        RECT  8.930 2.060 9.230 2.460 ;
        RECT  8.690 2.060 8.930 3.660 ;
        RECT  4.690 3.420 8.690 3.660 ;
        RECT  7.960 0.680 8.200 3.130 ;
        RECT  7.770 0.680 7.960 1.100 ;
        RECT  7.770 2.890 7.960 3.130 ;
        RECT  5.660 0.860 7.770 1.100 ;
        RECT  7.490 1.870 7.680 2.270 ;
        RECT  7.250 1.380 7.490 2.980 ;
        RECT  6.980 1.380 7.250 1.620 ;
        RECT  5.090 2.740 7.250 2.980 ;
        RECT  5.890 3.940 6.200 4.350 ;
        RECT  5.800 4.110 5.890 4.350 ;
        RECT  5.420 0.860 5.660 1.840 ;
        RECT  5.070 1.600 5.420 1.840 ;
        RECT  4.850 2.320 5.090 2.980 ;
        RECT  4.670 1.600 5.070 2.000 ;
        RECT  4.690 2.320 4.850 2.720 ;
        RECT  4.670 1.010 4.750 1.250 ;
        RECT  4.370 3.420 4.690 3.790 ;
        RECT  4.350 0.860 4.670 1.250 ;
        RECT  4.400 1.760 4.670 2.000 ;
        RECT  4.160 1.760 4.400 3.140 ;
        RECT  1.890 3.550 4.370 3.790 ;
        RECT  2.600 0.860 4.350 1.100 ;
        RECT  3.960 2.900 4.160 3.140 ;
        RECT  3.720 2.900 3.960 3.270 ;
        RECT  2.480 3.030 3.720 3.270 ;
        RECT  2.360 0.860 2.600 1.570 ;
        RECT  2.240 2.490 2.480 3.270 ;
        RECT  1.810 1.330 2.360 1.570 ;
        RECT  2.150 2.490 2.240 2.730 ;
        RECT  1.910 2.330 2.150 2.730 ;
        RECT  1.150 0.770 1.990 1.010 ;
        RECT  1.650 3.080 1.890 3.790 ;
        RECT  1.630 1.330 1.810 2.050 ;
        RECT  1.110 4.070 1.770 4.310 ;
        RECT  1.630 3.080 1.650 3.320 ;
        RECT  1.570 1.330 1.630 3.320 ;
        RECT  1.390 1.810 1.570 3.320 ;
        RECT  1.110 0.770 1.150 1.530 ;
        RECT  0.910 0.770 1.110 4.310 ;
        RECT  0.870 1.210 0.910 4.310 ;
    END
END TLATNSRX1

MACRO TLATNSXL
    CLASS CORE ;
    FOREIGN TLATNSXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.190 2.080 0.200 2.480 ;
        RECT  0.200 1.830 0.460 2.480 ;
        RECT  0.460 1.840 0.510 2.480 ;
        RECT  0.510 2.080 0.590 2.480 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  10.070 1.200 10.100 2.640 ;
        RECT  9.990 2.990 10.110 3.390 ;
        RECT  10.100 1.200 10.110 2.650 ;
        RECT  10.110 1.200 10.310 3.390 ;
        RECT  10.310 2.390 10.350 3.390 ;
        RECT  10.350 2.390 10.360 2.650 ;
        RECT  10.350 2.990 10.390 3.390 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  8.670 2.940 8.910 3.350 ;
        RECT  8.910 2.940 8.920 3.210 ;
        RECT  8.650 1.460 8.920 1.700 ;
        RECT  8.920 1.460 9.040 3.210 ;
        RECT  9.040 1.460 9.160 3.200 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  5.480 1.270 5.490 1.530 ;
        RECT  5.490 1.270 5.740 1.710 ;
        RECT  5.740 1.470 5.810 1.710 ;
        RECT  5.810 1.470 6.050 1.870 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.750 1.820 3.290 2.230 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.740 0.560 5.440 ;
        RECT  0.560 4.640 3.190 5.440 ;
        RECT  3.190 4.080 3.430 5.440 ;
        RECT  3.430 4.640 5.930 5.440 ;
        RECT  5.930 4.480 6.330 5.440 ;
        RECT  6.330 4.640 7.760 5.440 ;
        RECT  7.760 4.480 8.160 5.440 ;
        RECT  8.160 4.640 9.880 5.440 ;
        RECT  9.880 4.480 10.280 5.440 ;
        RECT  10.280 4.640 10.560 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 2.530 0.400 ;
        RECT  2.530 -0.400 2.930 0.560 ;
        RECT  2.930 -0.400 5.270 0.400 ;
        RECT  5.270 -0.400 5.670 0.560 ;
        RECT  5.670 -0.400 7.770 0.400 ;
        RECT  7.770 -0.400 8.170 0.560 ;
        RECT  8.170 -0.400 9.380 0.400 ;
        RECT  9.380 -0.400 9.780 0.560 ;
        RECT  9.780 -0.400 10.560 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  9.450 0.880 9.690 4.020 ;
        RECT  9.050 0.880 9.450 1.120 ;
        RECT  9.030 3.780 9.450 4.020 ;
        RECT  8.760 0.670 9.050 1.120 ;
        RECT  8.790 3.780 9.030 4.370 ;
        RECT  8.630 3.940 8.790 4.370 ;
        RECT  8.650 0.670 8.760 0.910 ;
        RECT  5.670 3.940 8.630 4.180 ;
        RECT  8.210 2.040 8.530 2.440 ;
        RECT  8.130 2.040 8.210 3.660 ;
        RECT  7.970 2.150 8.130 3.660 ;
        RECT  1.890 3.420 7.970 3.660 ;
        RECT  7.450 1.020 7.690 3.140 ;
        RECT  6.890 1.020 7.450 1.260 ;
        RECT  3.970 2.900 7.450 3.140 ;
        RECT  6.830 1.630 7.170 2.030 ;
        RECT  6.580 1.630 6.830 2.620 ;
        RECT  6.570 1.630 6.580 1.870 ;
        RECT  4.650 2.380 6.580 2.620 ;
        RECT  6.330 0.860 6.570 1.870 ;
        RECT  6.150 0.860 6.330 1.100 ;
        RECT  5.270 3.940 5.670 4.230 ;
        RECT  4.330 2.280 4.650 2.620 ;
        RECT  3.970 1.550 4.640 1.790 ;
        RECT  2.400 0.860 4.330 1.100 ;
        RECT  4.250 2.280 4.330 2.520 ;
        RECT  3.730 1.550 3.970 3.140 ;
        RECT  2.350 2.560 3.730 2.800 ;
        RECT  2.160 0.860 2.400 1.570 ;
        RECT  2.110 2.040 2.350 2.800 ;
        RECT  1.800 1.330 2.160 1.570 ;
        RECT  1.800 3.080 1.890 3.660 ;
        RECT  1.650 1.330 1.800 3.660 ;
        RECT  1.150 4.070 1.750 4.310 ;
        RECT  1.150 0.760 1.690 1.000 ;
        RECT  1.560 1.330 1.650 3.400 ;
        RECT  0.910 0.760 1.150 4.310 ;
    END
END TLATNSXL

MACRO TLATNSX4
    CLASS CORE ;
    FOREIGN TLATNSX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNSXL ;
    SIZE 14.520 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.210 2.650 ;
        RECT  0.210 2.060 0.460 2.650 ;
        RECT  0.460 2.060 0.540 2.640 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.650 1.820 12.850 3.220 ;
        RECT  12.850 1.390 13.000 3.220 ;
        RECT  13.000 1.230 13.090 3.250 ;
        RECT  13.090 2.850 13.400 3.250 ;
        RECT  13.090 1.230 13.400 1.630 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.330 1.820 11.450 3.220 ;
        RECT  11.450 1.400 11.460 3.220 ;
        RECT  11.460 1.230 11.780 3.250 ;
        RECT  11.780 2.850 11.860 3.250 ;
        RECT  11.780 1.230 11.860 1.630 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  6.800 1.270 6.810 1.530 ;
        RECT  6.810 1.270 7.060 1.710 ;
        RECT  7.060 1.470 7.500 1.710 ;
        RECT  7.500 1.470 7.740 1.870 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 1.830 2.980 2.090 ;
        RECT  2.980 1.830 2.990 2.300 ;
        RECT  2.990 1.830 3.390 2.530 ;
        RECT  3.390 1.830 3.400 2.300 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 3.270 5.440 ;
        RECT  3.270 3.940 3.670 5.440 ;
        RECT  3.670 4.640 7.640 5.440 ;
        RECT  7.640 4.480 8.040 5.440 ;
        RECT  8.040 4.640 9.380 5.440 ;
        RECT  9.380 4.480 9.780 5.440 ;
        RECT  9.780 4.640 10.730 5.440 ;
        RECT  10.730 4.480 11.130 5.440 ;
        RECT  11.130 4.640 12.270 5.440 ;
        RECT  12.270 4.210 12.670 5.440 ;
        RECT  12.670 4.640 13.670 5.440 ;
        RECT  13.670 4.210 14.070 5.440 ;
        RECT  14.070 4.640 14.520 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 2.360 0.400 ;
        RECT  2.360 -0.400 2.760 0.560 ;
        RECT  2.760 -0.400 4.940 0.400 ;
        RECT  4.940 -0.400 5.340 0.560 ;
        RECT  5.340 -0.400 7.080 0.400 ;
        RECT  7.080 -0.400 7.480 0.950 ;
        RECT  7.480 -0.400 9.350 0.400 ;
        RECT  9.350 -0.400 9.750 1.270 ;
        RECT  9.750 -0.400 10.850 0.400 ;
        RECT  10.850 -0.400 11.250 0.950 ;
        RECT  11.250 -0.400 12.270 0.400 ;
        RECT  12.270 -0.400 12.670 0.950 ;
        RECT  12.670 -0.400 13.670 0.400 ;
        RECT  13.670 -0.400 14.070 0.950 ;
        RECT  14.070 -0.400 14.520 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  13.640 2.200 13.880 3.920 ;
        RECT  13.570 2.200 13.640 2.440 ;
        RECT  10.600 3.680 13.640 3.920 ;
        RECT  13.330 2.040 13.570 2.440 ;
        RECT  10.820 1.350 11.060 3.050 ;
        RECT  10.510 1.350 10.820 1.590 ;
        RECT  10.600 2.810 10.820 3.050 ;
        RECT  10.440 2.810 10.600 3.930 ;
        RECT  10.140 2.040 10.540 2.440 ;
        RECT  10.110 1.190 10.510 1.590 ;
        RECT  10.200 2.810 10.440 4.180 ;
        RECT  7.360 3.940 10.200 4.180 ;
        RECT  9.870 2.200 10.140 2.440 ;
        RECT  9.630 2.200 9.870 3.660 ;
        RECT  1.850 3.420 9.630 3.660 ;
        RECT  9.070 2.900 9.170 3.140 ;
        RECT  8.830 0.950 9.070 3.140 ;
        RECT  8.590 0.950 8.830 1.190 ;
        RECT  5.980 2.900 8.830 3.140 ;
        RECT  8.430 1.600 8.550 2.000 ;
        RECT  8.310 1.600 8.430 2.620 ;
        RECT  8.070 0.860 8.310 2.620 ;
        RECT  7.840 0.860 8.070 1.100 ;
        RECT  8.060 1.840 8.070 2.620 ;
        RECT  6.660 2.380 8.060 2.620 ;
        RECT  6.960 3.940 7.360 4.250 ;
        RECT  6.260 2.280 6.660 2.620 ;
        RECT  5.980 1.500 6.390 1.740 ;
        RECT  5.210 0.860 6.120 1.100 ;
        RECT  5.740 1.500 5.980 3.140 ;
        RECT  4.250 2.670 5.740 2.910 ;
        RECT  4.970 0.860 5.210 1.250 ;
        RECT  2.480 1.010 4.970 1.250 ;
        RECT  4.010 2.670 4.250 3.050 ;
        RECT  2.500 2.810 4.010 3.050 ;
        RECT  2.260 2.370 2.500 3.050 ;
        RECT  2.240 1.010 2.480 1.570 ;
        RECT  2.110 2.370 2.260 2.610 ;
        RECT  1.750 1.330 2.240 1.570 ;
        RECT  1.870 2.210 2.110 2.610 ;
        RECT  1.170 0.760 1.960 1.000 ;
        RECT  1.610 2.890 1.850 3.660 ;
        RECT  1.590 1.330 1.750 1.930 ;
        RECT  1.590 2.890 1.610 3.130 ;
        RECT  1.510 1.330 1.590 3.130 ;
        RECT  1.350 1.690 1.510 3.130 ;
        RECT  1.060 3.510 1.190 3.750 ;
        RECT  1.060 0.760 1.170 1.410 ;
        RECT  0.930 0.760 1.060 3.750 ;
        RECT  0.820 1.170 0.930 3.750 ;
        RECT  0.770 1.170 0.820 1.410 ;
        RECT  0.790 3.510 0.820 3.750 ;
    END
END TLATNSX4

MACRO TLATNSX2
    CLASS CORE ;
    FOREIGN TLATNSX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNSXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.190 2.030 0.200 2.430 ;
        RECT  0.200 1.830 0.460 2.430 ;
        RECT  0.460 2.030 0.590 2.430 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  10.650 0.740 10.890 4.220 ;
        RECT  10.890 2.390 11.020 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.050 2.810 9.200 3.210 ;
        RECT  9.200 0.740 9.440 3.210 ;
        RECT  9.440 2.810 9.450 3.210 ;
        RECT  9.450 2.950 9.700 3.210 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  5.480 1.270 5.490 1.530 ;
        RECT  5.490 1.270 5.740 1.710 ;
        RECT  5.740 1.470 5.780 1.710 ;
        RECT  5.780 1.470 6.020 1.870 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 1.830 3.000 2.090 ;
        RECT  3.000 1.830 3.100 2.270 ;
        RECT  3.100 1.840 3.320 2.270 ;
        RECT  3.320 1.870 3.400 2.270 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.690 0.560 5.440 ;
        RECT  0.560 4.640 3.270 5.440 ;
        RECT  3.270 4.480 3.670 5.440 ;
        RECT  3.670 4.640 5.600 5.440 ;
        RECT  5.600 4.000 6.000 5.440 ;
        RECT  6.000 4.640 7.730 5.440 ;
        RECT  7.730 4.480 8.130 5.440 ;
        RECT  8.130 4.640 9.820 5.440 ;
        RECT  9.820 4.190 10.220 5.440 ;
        RECT  10.220 4.640 11.220 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 2.460 0.400 ;
        RECT  2.460 -0.400 2.860 0.560 ;
        RECT  2.860 -0.400 5.180 0.400 ;
        RECT  5.180 -0.400 5.580 0.560 ;
        RECT  5.580 -0.400 7.750 0.400 ;
        RECT  7.750 -0.400 7.990 1.350 ;
        RECT  7.990 -0.400 9.840 0.400 ;
        RECT  9.840 -0.400 10.240 1.580 ;
        RECT  10.240 -0.400 11.220 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.310 2.040 10.410 2.440 ;
        RECT  10.070 2.040 10.310 3.910 ;
        RECT  8.770 3.670 10.070 3.910 ;
        RECT  8.770 0.940 8.790 1.340 ;
        RECT  8.530 0.940 8.770 4.240 ;
        RECT  8.390 0.940 8.530 1.340 ;
        RECT  6.260 4.000 8.530 4.240 ;
        RECT  7.910 1.880 8.150 3.760 ;
        RECT  4.240 3.520 7.910 3.760 ;
        RECT  7.260 1.020 7.500 3.280 ;
        RECT  6.800 1.020 7.260 1.260 ;
        RECT  5.080 3.040 7.260 3.280 ;
        RECT  6.590 1.700 6.770 2.480 ;
        RECT  6.560 1.700 6.590 2.800 ;
        RECT  6.320 0.870 6.560 2.800 ;
        RECT  6.060 0.870 6.320 1.110 ;
        RECT  6.190 2.240 6.320 2.800 ;
        RECT  4.130 2.240 6.190 2.480 ;
        RECT  4.840 2.720 5.080 3.280 ;
        RECT  1.110 4.000 4.950 4.240 ;
        RECT  3.890 2.720 4.840 2.960 ;
        RECT  3.890 1.550 4.560 1.790 ;
        RECT  4.000 3.200 4.240 3.760 ;
        RECT  2.480 0.860 4.230 1.100 ;
        RECT  1.850 3.200 4.000 3.440 ;
        RECT  3.650 1.550 3.890 2.960 ;
        RECT  2.480 2.720 3.650 2.960 ;
        RECT  2.240 0.860 2.480 1.120 ;
        RECT  2.240 1.920 2.480 2.960 ;
        RECT  1.630 0.880 2.240 1.120 ;
        RECT  2.130 1.920 2.240 2.160 ;
        RECT  1.890 1.760 2.130 2.160 ;
        RECT  1.630 2.430 1.850 3.440 ;
        RECT  1.610 0.880 1.630 3.440 ;
        RECT  1.390 0.880 1.610 2.670 ;
        RECT  1.110 1.010 1.150 1.410 ;
        RECT  0.910 1.010 1.110 4.240 ;
        RECT  0.870 1.090 0.910 4.240 ;
    END
END TLATNSX2

MACRO TLATNSX1
    CLASS CORE ;
    FOREIGN TLATNSX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNSXL ;
    SIZE 9.900 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.190 1.950 0.200 2.490 ;
        RECT  0.200 1.830 0.460 2.490 ;
        RECT  0.460 2.090 0.590 2.490 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.330 1.300 9.350 1.700 ;
        RECT  9.340 2.990 9.450 3.390 ;
        RECT  9.440 2.390 9.450 2.650 ;
        RECT  9.350 1.300 9.450 1.820 ;
        RECT  9.450 1.300 9.690 3.390 ;
        RECT  9.690 2.390 9.700 2.650 ;
        RECT  9.690 1.300 9.730 1.950 ;
        RECT  9.690 2.990 9.740 3.390 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  7.690 1.480 7.890 1.720 ;
        RECT  7.890 1.480 8.110 3.200 ;
        RECT  8.110 1.480 8.130 3.430 ;
        RECT  8.130 2.940 8.350 3.430 ;
        RECT  8.350 2.940 8.370 3.210 ;
        RECT  8.370 2.950 8.380 3.210 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  5.240 2.020 5.480 2.500 ;
        RECT  5.480 2.260 5.730 2.650 ;
        RECT  5.730 2.390 5.740 2.650 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.660 1.960 2.740 2.360 ;
        RECT  2.740 1.840 2.840 2.360 ;
        RECT  2.840 1.830 3.060 2.360 ;
        RECT  3.060 1.830 3.100 2.090 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 3.100 5.440 ;
        RECT  3.100 4.200 3.500 5.440 ;
        RECT  3.500 4.640 5.530 5.440 ;
        RECT  5.530 4.480 5.930 5.440 ;
        RECT  5.930 4.640 8.750 5.440 ;
        RECT  8.750 4.480 9.150 5.440 ;
        RECT  9.150 4.640 9.900 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 2.280 0.400 ;
        RECT  2.280 -0.400 2.680 0.560 ;
        RECT  2.680 -0.400 4.860 0.400 ;
        RECT  4.860 -0.400 5.260 0.560 ;
        RECT  5.260 -0.400 6.900 0.400 ;
        RECT  6.900 -0.400 7.300 0.560 ;
        RECT  7.300 -0.400 8.740 0.400 ;
        RECT  8.740 -0.400 9.140 0.560 ;
        RECT  9.140 -0.400 9.900 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  8.740 0.800 8.980 3.940 ;
        RECT  8.160 0.800 8.740 1.040 ;
        RECT  8.430 3.700 8.740 3.940 ;
        RECT  8.190 3.700 8.430 4.360 ;
        RECT  8.030 4.120 8.190 4.360 ;
        RECT  7.760 0.680 8.160 1.040 ;
        RECT  4.740 0.800 7.760 1.040 ;
        RECT  7.360 2.260 7.600 4.370 ;
        RECT  6.410 4.130 7.360 4.370 ;
        RECT  7.050 1.280 7.120 3.760 ;
        RECT  6.880 1.280 7.050 3.840 ;
        RECT  6.240 1.280 6.880 1.520 ;
        RECT  6.650 3.520 6.880 3.840 ;
        RECT  4.670 3.520 6.650 3.760 ;
        RECT  6.440 1.780 6.640 3.110 ;
        RECT  6.400 1.780 6.440 3.280 ;
        RECT  6.170 4.000 6.410 4.370 ;
        RECT  6.000 1.780 6.400 2.020 ;
        RECT  6.120 2.870 6.400 3.280 ;
        RECT  4.140 4.000 6.170 4.240 ;
        RECT  5.150 3.040 6.120 3.280 ;
        RECT  5.760 1.280 6.000 2.020 ;
        RECT  5.520 1.280 5.760 1.520 ;
        RECT  4.910 2.750 5.150 3.280 ;
        RECT  4.050 2.750 4.910 2.990 ;
        RECT  4.610 0.800 4.740 2.310 ;
        RECT  4.430 3.230 4.670 3.760 ;
        RECT  4.500 0.800 4.610 2.390 ;
        RECT  4.370 1.990 4.500 2.390 ;
        RECT  3.730 3.230 4.430 3.470 ;
        RECT  3.730 1.360 4.260 1.600 ;
        RECT  3.900 3.710 4.140 4.240 ;
        RECT  2.560 0.800 3.930 1.040 ;
        RECT  1.890 3.710 3.900 3.950 ;
        RECT  3.490 1.360 3.730 3.470 ;
        RECT  2.420 3.230 3.490 3.470 ;
        RECT  2.320 0.800 2.560 1.500 ;
        RECT  2.190 2.490 2.420 3.470 ;
        RECT  1.670 1.260 2.320 1.500 ;
        RECT  2.180 1.960 2.190 3.470 ;
        RECT  1.950 1.960 2.180 2.730 ;
        RECT  1.150 0.690 2.040 0.930 ;
        RECT  1.670 3.080 1.890 3.950 ;
        RECT  1.650 1.260 1.670 3.950 ;
        RECT  1.430 1.260 1.650 3.400 ;
        RECT  1.150 4.120 1.410 4.360 ;
        RECT  0.910 0.690 1.150 4.360 ;
    END
END TLATNSX1

MACRO TLATNRXL
    CLASS CORE ;
    FOREIGN TLATNRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.250 2.390 3.490 3.390 ;
        RECT  3.490 2.390 3.510 2.640 ;
        RECT  3.510 2.390 4.160 2.630 ;
        RECT  4.160 2.390 4.240 2.650 ;
        RECT  4.240 1.880 4.420 2.650 ;
        RECT  4.420 1.880 4.480 2.630 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  7.330 1.220 7.370 1.620 ;
        RECT  7.370 1.220 7.460 1.820 ;
        RECT  7.310 3.160 7.470 3.560 ;
        RECT  7.460 1.220 7.470 2.090 ;
        RECT  7.470 1.220 7.710 3.560 ;
        RECT  7.710 1.220 7.720 2.090 ;
        RECT  7.720 1.220 7.730 1.960 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  5.910 0.670 5.990 0.910 ;
        RECT  6.050 3.480 6.290 4.170 ;
        RECT  5.990 0.670 6.310 1.100 ;
        RECT  6.290 3.480 6.400 3.770 ;
        RECT  6.400 3.480 6.780 3.720 ;
        RECT  6.310 0.860 6.780 1.100 ;
        RECT  6.780 0.860 7.020 3.720 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.180 1.830 0.600 2.520 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.980 2.240 2.440 2.660 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.530 5.440 ;
        RECT  1.530 3.840 1.930 5.440 ;
        RECT  1.930 4.640 3.570 5.440 ;
        RECT  3.570 4.110 3.970 5.440 ;
        RECT  3.970 4.640 5.180 5.440 ;
        RECT  5.180 4.480 5.580 5.440 ;
        RECT  5.580 4.640 6.720 5.440 ;
        RECT  6.720 4.480 7.120 5.440 ;
        RECT  7.120 4.640 7.920 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.780 0.400 ;
        RECT  1.780 -0.400 2.180 0.560 ;
        RECT  2.180 -0.400 5.190 0.400 ;
        RECT  5.190 -0.400 5.590 0.910 ;
        RECT  5.590 -0.400 6.700 0.400 ;
        RECT  6.700 -0.400 7.100 0.560 ;
        RECT  7.100 -0.400 7.920 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.280 1.470 6.520 3.180 ;
        RECT  5.980 1.470 6.280 1.710 ;
        RECT  5.970 2.780 6.280 3.180 ;
        RECT  5.470 2.940 5.970 3.180 ;
        RECT  5.520 2.040 5.920 2.440 ;
        RECT  4.990 2.120 5.520 2.360 ;
        RECT  5.230 2.940 5.470 3.910 ;
        RECT  4.820 3.670 5.230 3.910 ;
        RECT  4.750 1.180 4.990 3.290 ;
        RECT  3.760 1.180 4.750 1.420 ;
        RECT  4.310 3.050 4.750 3.290 ;
        RECT  4.150 3.050 4.310 3.450 ;
        RECT  3.910 3.050 4.150 3.870 ;
        RECT  3.110 3.630 3.910 3.870 ;
        RECT  3.480 1.660 3.880 2.050 ;
        RECT  3.440 0.980 3.760 1.420 ;
        RECT  3.010 1.660 3.480 1.900 ;
        RECT  3.360 0.980 3.440 1.220 ;
        RECT  2.790 3.630 3.110 4.160 ;
        RECT  2.770 1.660 3.010 3.310 ;
        RECT  2.710 3.760 2.790 4.160 ;
        RECT  1.810 1.660 2.770 1.900 ;
        RECT  2.440 3.070 2.770 3.310 ;
        RECT  1.740 0.870 1.810 1.900 ;
        RECT  1.500 0.870 1.740 3.540 ;
        RECT  1.310 0.870 1.500 1.130 ;
        RECT  1.060 3.300 1.500 3.540 ;
        RECT  0.910 0.770 1.310 1.130 ;
        RECT  1.190 2.180 1.260 2.580 ;
        RECT  1.150 2.180 1.190 3.040 ;
        RECT  0.950 1.410 1.150 3.040 ;
        RECT  0.820 3.300 1.060 4.080 ;
        RECT  0.910 1.410 0.950 2.420 ;
        RECT  0.790 2.800 0.950 3.040 ;
    END
END TLATNRXL

MACRO TLATNRX4
    CLASS CORE ;
    FOREIGN TLATNRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNRXL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.390 2.850 2.650 ;
        RECT  2.850 2.390 3.100 2.970 ;
        RECT  3.100 2.570 3.270 2.970 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  10.600 2.890 10.670 3.130 ;
        RECT  10.600 1.220 10.670 1.620 ;
        RECT  10.670 1.220 11.000 3.130 ;
        RECT  11.000 1.260 11.010 3.130 ;
        RECT  11.010 1.260 11.110 2.660 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.110 2.890 9.350 3.130 ;
        RECT  9.230 0.730 9.350 1.630 ;
        RECT  9.350 0.730 9.590 3.130 ;
        RECT  9.590 0.730 9.630 2.660 ;
        RECT  9.630 1.260 9.790 2.660 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  5.480 1.830 5.490 2.090 ;
        RECT  5.490 1.670 6.010 2.110 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.720 2.090 ;
        RECT  1.720 1.830 1.780 2.480 ;
        RECT  1.780 1.850 1.960 2.480 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 2.720 5.440 ;
        RECT  2.720 4.480 3.120 5.440 ;
        RECT  3.120 4.640 4.830 5.440 ;
        RECT  4.830 4.480 5.230 5.440 ;
        RECT  5.230 4.640 7.000 5.440 ;
        RECT  7.000 4.480 7.400 5.440 ;
        RECT  7.400 4.640 8.300 5.440 ;
        RECT  8.300 4.480 8.700 5.440 ;
        RECT  8.700 4.640 9.990 5.440 ;
        RECT  9.990 3.950 10.390 5.440 ;
        RECT  10.390 4.640 11.250 5.440 ;
        RECT  11.250 3.950 11.650 5.440 ;
        RECT  11.650 4.640 11.880 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.990 0.400 ;
        RECT  1.990 -0.400 2.390 1.010 ;
        RECT  2.390 -0.400 5.460 0.400 ;
        RECT  5.460 -0.400 6.540 0.560 ;
        RECT  6.540 -0.400 8.410 0.400 ;
        RECT  8.410 -0.400 8.810 0.560 ;
        RECT  8.810 -0.400 9.990 0.400 ;
        RECT  9.990 -0.400 10.390 0.940 ;
        RECT  10.390 -0.400 11.250 0.400 ;
        RECT  11.250 -0.400 11.650 0.940 ;
        RECT  11.650 -0.400 11.880 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  11.380 1.790 11.620 3.670 ;
        RECT  8.380 3.430 11.380 3.670 ;
        RECT  8.290 1.620 8.380 3.670 ;
        RECT  8.140 1.460 8.290 3.670 ;
        RECT  7.890 1.460 8.140 1.860 ;
        RECT  8.110 3.430 8.140 3.670 ;
        RECT  7.870 3.430 8.110 4.180 ;
        RECT  7.640 2.170 7.880 2.940 ;
        RECT  4.590 3.940 7.870 4.180 ;
        RECT  7.600 2.700 7.640 2.940 ;
        RECT  7.360 2.700 7.600 3.660 ;
        RECT  7.100 0.860 7.550 1.260 ;
        RECT  3.710 3.420 7.360 3.660 ;
        RECT  6.860 0.860 7.100 3.130 ;
        RECT  4.570 0.860 6.860 1.100 ;
        RECT  6.390 2.890 6.860 3.130 ;
        RECT  6.360 1.380 6.600 2.620 ;
        RECT  6.350 1.380 6.360 1.780 ;
        RECT  6.110 2.380 6.360 2.620 ;
        RECT  5.870 2.380 6.110 3.140 ;
        RECT  4.680 2.900 5.870 3.140 ;
        RECT  4.440 2.700 4.680 3.140 ;
        RECT  4.350 3.940 4.590 4.340 ;
        RECT  4.330 0.860 4.570 2.290 ;
        RECT  3.590 2.700 4.440 2.940 ;
        RECT  4.150 1.870 4.330 2.290 ;
        RECT  2.480 1.870 4.150 2.110 ;
        RECT  3.810 0.910 4.050 1.530 ;
        RECT  3.560 3.940 3.960 4.340 ;
        RECT  1.040 1.290 3.810 1.530 ;
        RECT  3.310 3.260 3.710 3.660 ;
        RECT  2.370 3.940 3.560 4.180 ;
        RECT  1.850 3.420 3.310 3.660 ;
        RECT  2.240 1.870 2.480 3.120 ;
        RECT  2.130 3.940 2.370 4.370 ;
        RECT  1.690 2.880 2.240 3.120 ;
        RECT  1.130 4.130 2.130 4.370 ;
        RECT  1.450 3.420 1.850 3.770 ;
        RECT  1.040 3.420 1.450 3.660 ;
        RECT  0.890 3.940 1.130 4.370 ;
        RECT  0.800 1.140 1.040 3.660 ;
        RECT  0.500 3.940 0.890 4.180 ;
        RECT  0.570 1.140 0.800 1.380 ;
        RECT  0.170 0.980 0.570 1.380 ;
        RECT  0.260 1.920 0.500 4.180 ;
    END
END TLATNRX4

MACRO TLATNRX2
    CLASS CORE ;
    FOREIGN TLATNRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNRXL ;
    SIZE 9.240 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.060 2.150 3.470 2.480 ;
        RECT  3.470 2.240 4.040 2.480 ;
        RECT  4.040 2.240 4.280 3.560 ;
        RECT  4.280 2.950 4.450 3.560 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  8.670 0.880 8.780 1.830 ;
        RECT  8.650 3.130 8.790 4.110 ;
        RECT  8.780 0.880 8.790 2.090 ;
        RECT  8.790 0.880 9.030 4.110 ;
        RECT  9.030 0.880 9.040 2.090 ;
        RECT  9.030 3.130 9.050 4.110 ;
        RECT  9.040 0.880 9.070 1.970 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  7.000 3.850 7.110 4.250 ;
        RECT  7.110 1.390 7.350 4.250 ;
        RECT  7.350 2.940 7.360 4.250 ;
        RECT  7.360 3.850 7.400 4.250 ;
        RECT  7.360 2.940 7.810 3.220 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.180 1.800 0.580 2.500 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 2.390 2.350 2.710 ;
        RECT  2.350 2.310 2.750 2.710 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.730 5.440 ;
        RECT  1.730 4.230 2.130 5.440 ;
        RECT  2.130 4.640 3.820 5.440 ;
        RECT  3.820 4.480 4.220 5.440 ;
        RECT  4.220 4.640 5.900 5.440 ;
        RECT  5.900 4.480 6.300 5.440 ;
        RECT  6.300 4.640 7.840 5.440 ;
        RECT  7.840 3.480 8.240 5.440 ;
        RECT  8.240 4.640 9.240 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 2.300 0.400 ;
        RECT  2.300 -0.400 2.700 0.560 ;
        RECT  2.700 -0.400 5.630 0.400 ;
        RECT  5.630 -0.400 6.030 0.560 ;
        RECT  6.030 -0.400 7.850 0.400 ;
        RECT  7.850 -0.400 8.250 0.560 ;
        RECT  8.250 -0.400 9.240 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  8.150 0.860 8.390 2.470 ;
        RECT  6.900 0.860 8.150 1.100 ;
        RECT  6.820 0.680 6.900 1.100 ;
        RECT  6.580 0.680 6.820 3.420 ;
        RECT  6.500 0.680 6.580 0.920 ;
        RECT  5.970 1.620 6.580 2.020 ;
        RECT  6.560 3.020 6.580 3.420 ;
        RECT  5.730 2.340 6.300 2.740 ;
        RECT  5.550 2.340 5.730 4.140 ;
        RECT  5.490 0.910 5.550 4.140 ;
        RECT  5.310 0.910 5.490 2.580 ;
        RECT  3.350 3.900 5.490 4.140 ;
        RECT  4.440 0.910 5.310 1.150 ;
        RECT  5.030 3.330 5.210 3.570 ;
        RECT  4.790 1.720 5.030 3.570 ;
        RECT  4.030 1.720 4.790 1.960 ;
        RECT  4.040 0.750 4.440 1.150 ;
        RECT  3.790 1.430 4.030 1.960 ;
        RECT  2.570 1.430 3.790 1.670 ;
        RECT  3.320 2.870 3.720 3.250 ;
        RECT  2.950 3.900 3.350 4.300 ;
        RECT  1.820 3.010 3.320 3.250 ;
        RECT  2.330 0.860 2.570 1.670 ;
        RECT  1.160 0.860 2.330 1.100 ;
        RECT  1.820 1.380 2.000 1.620 ;
        RECT  1.580 1.380 1.820 3.870 ;
        RECT  1.250 3.620 1.580 3.870 ;
        RECT  1.160 2.030 1.300 2.430 ;
        RECT  0.850 3.620 1.250 4.020 ;
        RECT  1.120 0.860 1.160 2.430 ;
        RECT  0.920 0.860 1.120 3.150 ;
        RECT  0.880 2.170 0.920 3.150 ;
    END
END TLATNRX2

MACRO TLATNRX1
    CLASS CORE ;
    FOREIGN TLATNRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNRXL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.250 2.390 3.490 3.360 ;
        RECT  3.490 2.390 3.510 2.640 ;
        RECT  3.510 2.390 4.160 2.630 ;
        RECT  4.160 2.390 4.240 2.650 ;
        RECT  4.240 1.860 4.420 2.650 ;
        RECT  4.420 1.860 4.480 2.630 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  7.330 1.170 7.460 1.570 ;
        RECT  7.310 2.930 7.470 3.330 ;
        RECT  7.460 1.170 7.470 2.090 ;
        RECT  7.470 1.170 7.710 3.330 ;
        RECT  7.710 1.170 7.720 2.090 ;
        RECT  7.720 1.170 7.730 1.570 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  5.910 0.670 5.990 0.910 ;
        RECT  6.050 3.480 6.290 4.170 ;
        RECT  5.990 0.670 6.310 1.100 ;
        RECT  6.290 3.480 6.400 3.770 ;
        RECT  6.400 3.480 6.780 3.720 ;
        RECT  6.310 0.860 6.780 1.100 ;
        RECT  6.780 0.860 7.020 3.720 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.180 1.830 0.600 2.520 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.980 2.270 2.450 2.660 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.530 5.440 ;
        RECT  1.530 3.760 1.930 5.440 ;
        RECT  1.930 4.640 3.570 5.440 ;
        RECT  3.570 4.110 3.970 5.440 ;
        RECT  3.970 4.640 5.180 5.440 ;
        RECT  5.180 4.480 5.580 5.440 ;
        RECT  5.580 4.640 6.720 5.440 ;
        RECT  6.720 4.480 7.120 5.440 ;
        RECT  7.120 4.640 7.920 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.780 0.400 ;
        RECT  1.780 -0.400 2.180 0.560 ;
        RECT  2.180 -0.400 5.190 0.400 ;
        RECT  5.190 -0.400 5.590 0.910 ;
        RECT  5.590 -0.400 6.700 0.400 ;
        RECT  6.700 -0.400 7.100 0.560 ;
        RECT  7.100 -0.400 7.920 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.280 1.470 6.520 3.180 ;
        RECT  5.980 1.470 6.280 1.710 ;
        RECT  5.970 2.780 6.280 3.180 ;
        RECT  5.470 2.940 5.970 3.180 ;
        RECT  5.520 2.040 5.920 2.440 ;
        RECT  4.990 2.120 5.520 2.360 ;
        RECT  5.230 2.940 5.470 3.910 ;
        RECT  4.820 3.670 5.230 3.910 ;
        RECT  4.750 1.180 4.990 3.290 ;
        RECT  3.760 1.180 4.750 1.420 ;
        RECT  4.310 3.050 4.750 3.290 ;
        RECT  4.150 3.050 4.310 3.450 ;
        RECT  3.910 3.050 4.150 3.860 ;
        RECT  3.110 3.620 3.910 3.860 ;
        RECT  3.480 1.660 3.880 2.050 ;
        RECT  3.440 0.980 3.760 1.420 ;
        RECT  3.010 1.660 3.480 1.900 ;
        RECT  3.360 0.980 3.440 1.220 ;
        RECT  2.790 3.620 3.110 4.130 ;
        RECT  2.770 1.660 3.010 3.210 ;
        RECT  2.710 3.730 2.790 4.130 ;
        RECT  1.810 1.660 2.770 1.900 ;
        RECT  2.440 2.970 2.770 3.210 ;
        RECT  1.740 0.870 1.810 1.900 ;
        RECT  1.500 0.870 1.740 3.520 ;
        RECT  1.310 0.870 1.500 1.110 ;
        RECT  1.130 3.280 1.500 3.520 ;
        RECT  0.910 0.770 1.310 1.110 ;
        RECT  1.150 2.180 1.260 3.040 ;
        RECT  1.020 1.410 1.150 3.040 ;
        RECT  0.890 3.280 1.130 4.060 ;
        RECT  0.910 1.410 1.020 2.420 ;
        RECT  0.790 2.800 1.020 3.040 ;
    END
END TLATNRX1

MACRO TLATNXL
    CLASS CORE ;
    FOREIGN TLATNXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.670 1.140 6.800 1.540 ;
        RECT  6.680 3.060 6.810 3.460 ;
        RECT  6.800 1.140 6.810 2.090 ;
        RECT  6.810 1.140 7.050 3.460 ;
        RECT  7.050 1.140 7.060 2.090 ;
        RECT  7.060 1.140 7.070 1.540 ;
        RECT  7.050 3.060 7.080 3.460 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  5.070 0.690 5.470 1.100 ;
        RECT  5.470 0.720 5.490 1.100 ;
        RECT  5.340 3.480 5.580 4.180 ;
        RECT  5.580 3.480 5.740 3.770 ;
        RECT  5.740 3.480 6.140 3.720 ;
        RECT  5.490 0.860 6.140 1.100 ;
        RECT  6.140 0.860 6.380 3.720 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.460 2.520 ;
        RECT  0.460 1.900 0.610 2.520 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.090 2.060 2.490 2.650 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.740 0.560 5.440 ;
        RECT  0.560 4.640 1.790 5.440 ;
        RECT  1.790 4.110 2.190 5.440 ;
        RECT  2.190 4.640 4.450 5.440 ;
        RECT  4.450 4.480 4.850 5.440 ;
        RECT  4.850 4.640 6.050 5.440 ;
        RECT  6.050 4.480 6.450 5.440 ;
        RECT  6.450 4.640 7.260 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.780 0.400 ;
        RECT  1.780 -0.400 2.180 0.560 ;
        RECT  2.180 -0.400 4.200 0.400 ;
        RECT  4.200 -0.400 4.600 0.560 ;
        RECT  4.600 -0.400 5.980 0.400 ;
        RECT  5.980 -0.400 6.380 0.560 ;
        RECT  6.380 -0.400 7.260 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.720 2.070 5.860 2.470 ;
        RECT  5.700 2.070 5.720 3.210 ;
        RECT  5.460 1.460 5.700 3.210 ;
        RECT  5.070 1.460 5.460 1.700 ;
        RECT  5.320 2.810 5.460 3.210 ;
        RECT  4.990 2.970 5.320 3.210 ;
        RECT  4.470 2.040 5.140 2.440 ;
        RECT  4.750 2.970 4.990 4.060 ;
        RECT  4.090 3.820 4.750 4.060 ;
        RECT  4.230 0.880 4.470 3.540 ;
        RECT  3.070 0.880 4.230 1.120 ;
        RECT  3.390 3.300 4.230 3.540 ;
        RECT  3.480 1.550 3.770 1.790 ;
        RECT  3.240 1.550 3.480 2.960 ;
        RECT  3.150 3.300 3.390 3.800 ;
        RECT  1.810 1.550 3.240 1.790 ;
        RECT  2.810 2.720 3.240 2.960 ;
        RECT  1.670 0.860 1.810 2.950 ;
        RECT  1.570 0.860 1.670 3.840 ;
        RECT  1.310 0.860 1.570 1.100 ;
        RECT  1.430 2.710 1.570 3.840 ;
        RECT  1.310 3.600 1.430 3.840 ;
        RECT  0.990 0.680 1.310 1.100 ;
        RECT  0.910 3.600 1.310 4.000 ;
        RECT  1.150 2.030 1.290 2.430 ;
        RECT  0.910 1.380 1.150 3.170 ;
        RECT  0.910 0.680 0.990 0.920 ;
    END
END TLATNXL

MACRO TLATNX4
    CLASS CORE ;
    FOREIGN TLATNX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.840 1.370 10.000 1.770 ;
        RECT  10.000 1.370 10.240 3.270 ;
        RECT  10.240 1.530 10.450 3.270 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  8.510 2.870 8.690 3.270 ;
        RECT  8.460 1.450 8.690 1.690 ;
        RECT  8.690 1.450 8.910 3.270 ;
        RECT  8.910 1.450 9.030 3.220 ;
        RECT  9.030 1.820 9.130 3.220 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.160 1.860 0.200 2.530 ;
        RECT  0.200 1.860 0.460 2.650 ;
        RECT  0.460 1.860 0.490 2.640 ;
        RECT  0.490 1.860 0.570 2.530 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.410 2.330 4.070 2.570 ;
        RECT  4.070 1.960 4.160 2.570 ;
        RECT  4.160 1.960 4.260 2.650 ;
        RECT  4.260 1.960 4.360 3.030 ;
        RECT  4.360 1.690 4.600 3.030 ;
        RECT  4.600 2.790 4.680 3.030 ;
        RECT  4.600 1.690 4.980 1.930 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.870 5.440 ;
        RECT  1.870 4.240 2.270 5.440 ;
        RECT  2.270 4.640 4.230 5.440 ;
        RECT  4.230 4.230 4.630 5.440 ;
        RECT  4.630 4.640 6.660 5.440 ;
        RECT  6.660 4.480 7.060 5.440 ;
        RECT  7.060 4.640 7.770 5.440 ;
        RECT  7.770 4.480 8.170 5.440 ;
        RECT  8.170 4.640 9.280 5.440 ;
        RECT  9.280 4.130 9.680 5.440 ;
        RECT  9.680 4.640 10.640 5.440 ;
        RECT  10.640 4.130 11.040 5.440 ;
        RECT  11.040 4.640 11.220 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 2.090 0.400 ;
        RECT  2.090 -0.400 2.490 0.560 ;
        RECT  2.490 -0.400 4.520 0.400 ;
        RECT  4.520 -0.400 4.920 0.970 ;
        RECT  4.920 -0.400 7.020 0.400 ;
        RECT  7.020 -0.400 7.420 0.560 ;
        RECT  7.420 -0.400 9.130 0.400 ;
        RECT  9.130 -0.400 9.530 1.090 ;
        RECT  9.530 -0.400 10.560 0.400 ;
        RECT  10.560 -0.400 10.960 1.090 ;
        RECT  10.960 -0.400 11.220 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.690 2.250 10.930 3.850 ;
        RECT  8.040 3.610 10.690 3.850 ;
        RECT  7.800 1.540 8.040 3.850 ;
        RECT  7.490 1.540 7.800 1.780 ;
        RECT  6.970 2.860 7.800 3.260 ;
        RECT  6.690 2.320 7.540 2.560 ;
        RECT  7.090 1.380 7.490 1.780 ;
        RECT  6.320 3.020 6.970 3.260 ;
        RECT  6.450 1.050 6.690 2.560 ;
        RECT  5.620 1.050 6.450 1.290 ;
        RECT  5.980 2.320 6.450 2.560 ;
        RECT  5.970 1.610 6.210 2.010 ;
        RECT  5.740 2.320 5.980 3.990 ;
        RECT  5.500 1.770 5.970 2.010 ;
        RECT  3.450 3.750 5.740 3.990 ;
        RECT  5.380 1.050 5.620 1.450 ;
        RECT  5.260 1.770 5.500 3.240 ;
        RECT  3.740 1.210 5.380 1.450 ;
        RECT  5.160 3.000 5.260 3.240 ;
        RECT  4.920 3.000 5.160 3.510 ;
        RECT  3.980 3.270 4.920 3.510 ;
        RECT  3.740 2.930 3.980 3.510 ;
        RECT  3.340 1.090 3.740 1.450 ;
        RECT  2.860 1.850 3.740 2.090 ;
        RECT  3.680 2.930 3.740 3.170 ;
        RECT  3.360 2.920 3.680 3.170 ;
        RECT  3.050 3.440 3.450 4.340 ;
        RECT  1.850 2.920 3.360 3.160 ;
        RECT  2.620 0.910 2.860 2.090 ;
        RECT  1.070 0.910 2.620 1.150 ;
        RECT  1.850 1.450 1.900 1.690 ;
        RECT  1.610 1.450 1.850 3.250 ;
        RECT  1.500 1.450 1.610 1.690 ;
        RECT  1.370 2.840 1.610 3.250 ;
        RECT  1.070 1.930 1.260 2.330 ;
        RECT  0.830 0.910 1.070 3.990 ;
    END
END TLATNX4

MACRO TLATNX2
    CLASS CORE ;
    FOREIGN TLATNX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNXL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  8.010 1.170 8.120 1.570 ;
        RECT  7.800 3.130 8.130 4.110 ;
        RECT  8.120 1.170 8.130 2.090 ;
        RECT  8.130 1.170 8.200 4.110 ;
        RECT  8.200 1.170 8.370 4.100 ;
        RECT  8.370 1.170 8.380 2.090 ;
        RECT  8.380 1.170 8.410 1.570 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.080 3.760 6.370 4.250 ;
        RECT  6.370 1.380 6.610 4.250 ;
        RECT  6.610 2.940 7.060 3.220 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.210 2.090 ;
        RECT  0.210 1.800 0.610 2.520 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 2.390 2.190 2.650 ;
        RECT  2.190 2.390 2.360 2.710 ;
        RECT  2.360 2.300 2.680 2.710 ;
        RECT  2.680 2.300 2.760 2.700 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.740 0.560 5.440 ;
        RECT  0.560 4.640 2.180 5.440 ;
        RECT  2.180 4.150 2.580 5.440 ;
        RECT  2.580 4.640 4.930 5.440 ;
        RECT  4.930 4.480 5.330 5.440 ;
        RECT  5.330 4.640 6.960 5.440 ;
        RECT  6.960 3.480 7.360 5.440 ;
        RECT  7.360 4.640 8.580 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 2.290 0.400 ;
        RECT  2.290 -0.400 2.690 0.560 ;
        RECT  2.690 -0.400 4.710 0.400 ;
        RECT  4.710 -0.400 5.110 0.560 ;
        RECT  5.110 -0.400 7.160 0.400 ;
        RECT  7.160 -0.400 7.560 0.560 ;
        RECT  7.560 -0.400 8.580 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  7.390 2.070 7.760 2.470 ;
        RECT  7.360 0.860 7.390 2.470 ;
        RECT  7.150 0.860 7.360 2.390 ;
        RECT  5.980 0.860 7.150 1.100 ;
        RECT  5.880 0.680 5.980 1.100 ;
        RECT  5.640 0.680 5.880 3.310 ;
        RECT  5.580 0.680 5.640 0.920 ;
        RECT  5.370 1.600 5.640 2.000 ;
        RECT  5.090 2.320 5.360 2.720 ;
        RECT  4.850 0.910 5.090 4.020 ;
        RECT  3.980 0.910 4.850 1.150 ;
        RECT  3.920 3.780 4.850 4.020 ;
        RECT  4.330 1.900 4.570 3.500 ;
        RECT  3.720 1.900 4.330 2.140 ;
        RECT  3.860 3.260 4.330 3.500 ;
        RECT  3.810 2.460 4.050 2.860 ;
        RECT  3.580 0.750 3.980 1.150 ;
        RECT  3.520 3.780 3.920 4.220 ;
        RECT  3.370 2.620 3.810 2.860 ;
        RECT  3.560 1.740 3.720 2.140 ;
        RECT  3.320 1.430 3.560 2.140 ;
        RECT  3.130 2.620 3.370 3.250 ;
        RECT  2.580 1.430 3.320 1.670 ;
        RECT  1.820 3.010 3.130 3.250 ;
        RECT  2.340 0.860 2.580 1.670 ;
        RECT  1.160 0.860 2.340 1.100 ;
        RECT  1.820 1.380 2.060 1.620 ;
        RECT  1.580 1.380 1.820 4.070 ;
        RECT  1.350 3.670 1.580 4.070 ;
        RECT  1.160 2.030 1.290 2.430 ;
        RECT  0.920 0.860 1.160 3.150 ;
        RECT  0.850 2.750 0.920 3.150 ;
    END
END TLATNX2

MACRO TLATNX1
    CLASS CORE ;
    FOREIGN TLATNX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATNXL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.690 1.170 6.800 1.850 ;
        RECT  6.690 2.930 6.810 3.330 ;
        RECT  6.800 1.170 6.810 2.090 ;
        RECT  6.810 1.170 7.050 3.330 ;
        RECT  7.050 1.170 7.060 2.090 ;
        RECT  7.050 2.930 7.090 3.330 ;
        RECT  7.060 1.170 7.090 1.570 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  5.320 3.770 5.400 4.170 ;
        RECT  5.180 0.670 5.470 0.910 ;
        RECT  5.400 3.520 5.480 4.170 ;
        RECT  5.470 0.670 5.710 1.100 ;
        RECT  5.480 3.510 5.720 4.170 ;
        RECT  5.720 3.510 5.740 3.770 ;
        RECT  5.740 3.520 6.170 3.760 ;
        RECT  5.710 0.860 6.170 1.100 ;
        RECT  6.170 0.860 6.410 3.760 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.180 1.960 0.200 2.520 ;
        RECT  0.200 1.830 0.460 2.520 ;
        RECT  0.460 1.960 0.580 2.520 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.150 2.570 2.180 2.970 ;
        RECT  2.180 2.390 2.440 2.970 ;
        RECT  2.440 2.570 2.550 2.970 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.770 0.560 5.440 ;
        RECT  0.560 4.640 1.910 5.440 ;
        RECT  1.910 3.720 2.310 5.440 ;
        RECT  2.310 4.640 4.510 5.440 ;
        RECT  4.510 4.480 4.910 5.440 ;
        RECT  4.910 4.640 6.080 5.440 ;
        RECT  6.080 4.480 6.480 5.440 ;
        RECT  6.480 4.640 7.260 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.840 0.400 ;
        RECT  1.840 -0.400 2.240 0.560 ;
        RECT  2.240 -0.400 4.310 0.400 ;
        RECT  4.310 -0.400 4.710 0.560 ;
        RECT  4.710 -0.400 5.980 0.400 ;
        RECT  5.980 -0.400 6.380 0.560 ;
        RECT  6.380 -0.400 7.260 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.650 1.470 5.890 3.190 ;
        RECT  5.200 1.470 5.650 1.710 ;
        RECT  5.320 2.780 5.650 3.190 ;
        RECT  4.960 2.950 5.320 3.190 ;
        RECT  4.440 2.040 5.250 2.440 ;
        RECT  4.720 2.950 4.960 4.110 ;
        RECT  4.150 3.870 4.720 4.110 ;
        RECT  4.200 0.860 4.440 3.510 ;
        RECT  3.530 0.860 4.200 1.100 ;
        RECT  3.530 3.270 4.200 3.510 ;
        RECT  3.670 1.470 3.840 1.870 ;
        RECT  3.430 1.470 3.670 2.950 ;
        RECT  3.130 0.700 3.530 1.100 ;
        RECT  3.130 3.270 3.530 3.670 ;
        RECT  1.810 1.470 3.430 1.710 ;
        RECT  2.870 2.710 3.430 2.950 ;
        RECT  1.630 0.870 1.810 3.170 ;
        RECT  1.570 0.870 1.630 4.120 ;
        RECT  1.370 0.870 1.570 1.110 ;
        RECT  1.390 2.930 1.570 4.120 ;
        RECT  1.100 3.720 1.390 4.120 ;
        RECT  0.970 0.740 1.370 1.110 ;
        RECT  1.150 2.240 1.290 2.640 ;
        RECT  1.110 1.380 1.150 2.640 ;
        RECT  0.910 1.380 1.110 3.320 ;
        RECT  0.870 2.320 0.910 3.320 ;
    END
END TLATNX1

MACRO TLATXL
    CLASS CORE ;
    FOREIGN TLATXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.650 3.060 6.810 3.460 ;
        RECT  6.800 1.830 6.810 2.090 ;
        RECT  6.690 1.140 6.810 1.540 ;
        RECT  6.810 1.140 7.050 3.460 ;
        RECT  7.050 1.830 7.060 2.090 ;
        RECT  7.050 1.140 7.090 1.540 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  5.100 3.780 5.260 4.180 ;
        RECT  5.160 0.690 5.470 0.930 ;
        RECT  5.260 3.540 5.480 4.180 ;
        RECT  5.480 3.510 5.500 4.180 ;
        RECT  5.500 3.510 5.590 3.780 ;
        RECT  5.470 0.690 5.710 1.040 ;
        RECT  5.590 3.500 5.720 3.780 ;
        RECT  5.720 3.500 5.740 3.770 ;
        RECT  5.740 3.500 5.830 3.760 ;
        RECT  5.830 3.500 5.920 3.740 ;
        RECT  5.710 0.800 5.920 1.040 ;
        RECT  5.920 0.800 6.160 3.740 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.460 2.620 ;
        RECT  0.460 1.840 0.600 2.620 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.080 2.320 2.600 2.860 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.690 0.560 5.440 ;
        RECT  0.560 4.640 1.790 5.440 ;
        RECT  1.790 4.120 2.190 5.440 ;
        RECT  2.190 4.640 4.290 5.440 ;
        RECT  4.290 4.480 4.690 5.440 ;
        RECT  4.690 4.640 6.020 5.440 ;
        RECT  6.020 4.480 6.420 5.440 ;
        RECT  6.420 4.640 7.260 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.790 0.400 ;
        RECT  1.790 -0.400 2.190 0.560 ;
        RECT  2.190 -0.400 4.290 0.400 ;
        RECT  4.290 -0.400 4.690 0.560 ;
        RECT  4.690 -0.400 5.980 0.400 ;
        RECT  5.980 -0.400 6.380 0.560 ;
        RECT  6.380 -0.400 7.260 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.440 1.460 5.680 3.160 ;
        RECT  5.160 1.460 5.440 1.700 ;
        RECT  4.710 2.920 5.440 3.160 ;
        RECT  4.640 2.010 5.040 2.440 ;
        RECT  4.470 2.920 4.710 3.830 ;
        RECT  4.190 2.010 4.640 2.270 ;
        RECT  4.330 3.590 4.470 3.830 ;
        RECT  3.930 3.590 4.330 3.990 ;
        RECT  3.950 2.010 4.190 3.290 ;
        RECT  3.820 2.010 3.950 2.250 ;
        RECT  3.530 3.050 3.950 3.290 ;
        RECT  3.580 0.670 3.820 2.250 ;
        RECT  3.300 2.530 3.670 2.770 ;
        RECT  3.140 0.670 3.580 0.910 ;
        RECT  3.290 3.050 3.530 4.190 ;
        RECT  3.210 1.320 3.300 2.770 ;
        RECT  3.130 3.790 3.290 4.190 ;
        RECT  3.060 1.240 3.210 2.770 ;
        RECT  2.810 1.240 3.060 1.640 ;
        RECT  1.810 1.390 2.810 1.630 ;
        RECT  1.670 0.860 1.810 3.140 ;
        RECT  1.570 0.860 1.670 3.840 ;
        RECT  1.310 0.860 1.570 1.100 ;
        RECT  1.430 2.900 1.570 3.840 ;
        RECT  1.310 3.600 1.430 3.840 ;
        RECT  0.910 0.680 1.310 1.100 ;
        RECT  0.910 3.600 1.310 4.000 ;
        RECT  1.150 2.030 1.290 2.430 ;
        RECT  0.910 1.380 1.150 3.170 ;
    END
END TLATXL

MACRO TLATX4
    CLASS CORE ;
    FOREIGN TLATX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.840 1.370 10.000 1.770 ;
        RECT  10.000 1.370 10.240 3.270 ;
        RECT  10.240 1.530 10.450 3.270 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  8.510 2.870 8.690 3.270 ;
        RECT  8.460 1.450 8.690 1.690 ;
        RECT  8.690 1.450 8.910 3.270 ;
        RECT  8.910 1.450 9.030 3.220 ;
        RECT  9.030 1.820 9.130 3.220 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.130 1.860 0.460 2.650 ;
        RECT  0.460 1.860 0.490 2.640 ;
        RECT  0.490 1.860 0.570 2.530 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.410 2.330 4.070 2.570 ;
        RECT  4.070 1.960 4.160 2.570 ;
        RECT  4.160 1.960 4.260 2.650 ;
        RECT  4.260 1.960 4.360 3.030 ;
        RECT  4.360 1.690 4.600 3.030 ;
        RECT  4.600 2.790 4.680 3.030 ;
        RECT  4.600 1.690 4.980 1.930 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.870 5.440 ;
        RECT  1.870 4.240 2.270 5.440 ;
        RECT  2.270 4.640 4.230 5.440 ;
        RECT  4.230 4.230 4.630 5.440 ;
        RECT  4.630 4.640 6.660 5.440 ;
        RECT  6.660 4.480 7.060 5.440 ;
        RECT  7.060 4.640 7.770 5.440 ;
        RECT  7.770 4.480 8.170 5.440 ;
        RECT  8.170 4.640 9.280 5.440 ;
        RECT  9.280 4.130 9.680 5.440 ;
        RECT  9.680 4.640 10.640 5.440 ;
        RECT  10.640 4.130 11.040 5.440 ;
        RECT  11.040 4.640 11.220 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 2.090 0.400 ;
        RECT  2.090 -0.400 2.490 0.560 ;
        RECT  2.490 -0.400 4.520 0.400 ;
        RECT  4.520 -0.400 4.920 0.970 ;
        RECT  4.920 -0.400 7.020 0.400 ;
        RECT  7.020 -0.400 7.420 0.560 ;
        RECT  7.420 -0.400 9.130 0.400 ;
        RECT  9.130 -0.400 9.530 1.090 ;
        RECT  9.530 -0.400 10.560 0.400 ;
        RECT  10.560 -0.400 10.960 1.090 ;
        RECT  10.960 -0.400 11.220 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.690 2.250 10.930 3.850 ;
        RECT  8.040 3.610 10.690 3.850 ;
        RECT  7.800 1.540 8.040 3.850 ;
        RECT  7.490 1.540 7.800 1.780 ;
        RECT  6.970 2.860 7.800 3.260 ;
        RECT  6.690 2.320 7.540 2.560 ;
        RECT  7.090 1.380 7.490 1.780 ;
        RECT  6.320 3.020 6.970 3.260 ;
        RECT  6.450 1.050 6.690 2.560 ;
        RECT  5.620 1.050 6.450 1.290 ;
        RECT  5.980 2.320 6.450 2.560 ;
        RECT  5.970 1.610 6.210 2.010 ;
        RECT  5.740 2.320 5.980 3.990 ;
        RECT  5.500 1.770 5.970 2.010 ;
        RECT  3.450 3.750 5.740 3.990 ;
        RECT  5.380 1.050 5.620 1.450 ;
        RECT  5.260 1.770 5.500 3.240 ;
        RECT  3.740 1.210 5.380 1.450 ;
        RECT  5.160 3.000 5.260 3.240 ;
        RECT  4.920 3.000 5.160 3.510 ;
        RECT  3.980 3.270 4.920 3.510 ;
        RECT  3.740 2.930 3.980 3.510 ;
        RECT  3.340 1.090 3.740 1.450 ;
        RECT  1.850 1.850 3.740 2.090 ;
        RECT  3.680 2.930 3.740 3.170 ;
        RECT  3.360 2.920 3.680 3.170 ;
        RECT  3.050 3.440 3.450 4.340 ;
        RECT  2.460 2.920 3.360 3.160 ;
        RECT  2.220 2.920 2.460 3.910 ;
        RECT  1.070 3.670 2.220 3.910 ;
        RECT  1.610 1.370 1.850 3.250 ;
        RECT  1.580 1.370 1.610 1.770 ;
        RECT  1.370 2.840 1.610 3.250 ;
        RECT  1.070 1.930 1.260 2.330 ;
        RECT  0.830 1.290 1.070 3.990 ;
    END
END TLATX4

MACRO TLATX2
    CLASS CORE ;
    FOREIGN TLATX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATXL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  7.860 0.810 8.030 1.790 ;
        RECT  8.030 0.810 8.120 1.820 ;
        RECT  7.860 3.120 8.130 4.100 ;
        RECT  8.120 0.810 8.130 2.090 ;
        RECT  8.130 0.810 8.260 4.100 ;
        RECT  8.260 0.810 8.370 4.090 ;
        RECT  8.370 1.830 8.380 2.090 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.140 3.850 6.220 4.330 ;
        RECT  6.220 1.390 6.460 4.330 ;
        RECT  6.460 3.850 6.540 4.330 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.170 2.020 0.200 2.620 ;
        RECT  0.200 1.830 0.460 2.620 ;
        RECT  0.460 2.020 0.570 2.620 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 2.390 2.190 2.650 ;
        RECT  2.190 2.390 2.500 2.700 ;
        RECT  2.500 2.300 2.900 2.700 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.730 0.560 5.440 ;
        RECT  0.560 4.640 2.260 5.440 ;
        RECT  2.260 4.050 2.660 5.440 ;
        RECT  2.660 4.640 5.040 5.440 ;
        RECT  5.040 4.480 5.440 5.440 ;
        RECT  5.440 4.640 7.020 5.440 ;
        RECT  7.020 3.480 7.420 5.440 ;
        RECT  7.420 4.640 8.580 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 2.250 0.400 ;
        RECT  2.250 -0.400 2.650 0.560 ;
        RECT  2.650 -0.400 4.730 0.400 ;
        RECT  4.730 -0.400 5.130 0.560 ;
        RECT  5.130 -0.400 7.020 0.400 ;
        RECT  7.020 -0.400 7.420 0.560 ;
        RECT  7.420 -0.400 8.580 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  7.450 2.070 7.610 2.470 ;
        RECT  7.210 0.860 7.450 2.470 ;
        RECT  6.020 0.860 7.210 1.100 ;
        RECT  5.940 0.680 6.020 1.100 ;
        RECT  5.700 0.680 5.940 3.310 ;
        RECT  5.620 0.680 5.700 0.920 ;
        RECT  5.040 1.600 5.700 2.000 ;
        RECT  4.730 2.320 5.420 2.720 ;
        RECT  4.490 0.910 4.730 4.300 ;
        RECT  3.580 0.910 4.490 1.150 ;
        RECT  3.500 4.060 4.490 4.300 ;
        RECT  3.660 3.470 4.210 3.710 ;
        RECT  3.940 1.430 4.180 2.990 ;
        RECT  2.560 1.430 3.940 1.670 ;
        RECT  3.420 1.950 3.660 3.710 ;
        RECT  3.260 1.950 3.420 2.190 ;
        RECT  1.820 3.470 3.420 3.710 ;
        RECT  2.320 0.860 2.560 1.670 ;
        RECT  1.150 0.860 2.320 1.100 ;
        RECT  1.820 1.380 1.980 1.620 ;
        RECT  1.580 1.380 1.820 4.080 ;
        RECT  1.380 3.680 1.580 4.080 ;
        RECT  1.150 2.030 1.290 2.430 ;
        RECT  0.910 0.860 1.150 3.150 ;
        RECT  0.860 2.750 0.910 3.150 ;
    END
END TLATX2

MACRO TLATX1
    CLASS CORE ;
    FOREIGN TLATX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TLATXL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.670 1.170 6.800 1.570 ;
        RECT  6.670 2.930 6.810 3.330 ;
        RECT  6.800 1.170 6.810 2.090 ;
        RECT  6.810 1.170 7.050 3.330 ;
        RECT  7.050 1.170 7.060 2.090 ;
        RECT  7.050 2.930 7.070 3.330 ;
        RECT  7.060 1.170 7.070 1.570 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  5.210 3.770 5.370 4.170 ;
        RECT  5.150 0.680 5.420 0.920 ;
        RECT  5.370 3.520 5.480 4.170 ;
        RECT  5.480 3.510 5.610 4.170 ;
        RECT  5.420 0.680 5.660 1.100 ;
        RECT  5.610 3.510 5.740 3.770 ;
        RECT  5.740 3.520 6.150 3.760 ;
        RECT  5.660 0.860 6.150 1.100 ;
        RECT  6.150 0.860 6.390 3.760 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.210 2.090 ;
        RECT  0.210 1.830 0.460 2.620 ;
        RECT  0.460 2.010 0.630 2.620 ;
        RECT  0.630 2.310 0.640 2.620 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 2.390 2.190 2.650 ;
        RECT  2.190 2.390 2.440 2.960 ;
        RECT  2.440 2.560 2.600 2.960 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.960 5.440 ;
        RECT  1.960 3.710 2.360 5.440 ;
        RECT  2.360 4.640 4.400 5.440 ;
        RECT  4.400 4.480 4.800 5.440 ;
        RECT  4.800 4.640 6.040 5.440 ;
        RECT  6.040 4.480 6.440 5.440 ;
        RECT  6.440 4.640 7.260 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.800 0.400 ;
        RECT  1.800 -0.400 2.200 0.560 ;
        RECT  2.200 -0.400 4.330 0.400 ;
        RECT  4.330 -0.400 4.730 0.560 ;
        RECT  4.730 -0.400 5.970 0.400 ;
        RECT  5.970 -0.400 6.370 0.560 ;
        RECT  6.370 -0.400 7.260 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.490 1.470 5.730 3.200 ;
        RECT  5.210 1.470 5.490 1.710 ;
        RECT  5.210 2.800 5.490 3.200 ;
        RECT  4.820 2.960 5.210 3.200 ;
        RECT  4.300 2.040 5.090 2.440 ;
        RECT  4.580 2.960 4.820 3.980 ;
        RECT  4.040 3.740 4.580 3.980 ;
        RECT  4.060 2.040 4.300 3.460 ;
        RECT  3.940 2.040 4.060 2.280 ;
        RECT  3.630 3.220 4.060 3.460 ;
        RECT  3.700 0.850 3.940 2.280 ;
        RECT  3.220 2.640 3.780 2.880 ;
        RECT  3.570 0.850 3.700 1.090 ;
        RECT  3.390 3.220 3.630 4.370 ;
        RECT  3.170 0.690 3.570 1.090 ;
        RECT  3.230 3.970 3.390 4.370 ;
        RECT  2.980 1.400 3.220 2.880 ;
        RECT  2.820 1.400 2.980 1.800 ;
        RECT  1.810 1.480 2.820 1.720 ;
        RECT  1.670 0.870 1.810 3.160 ;
        RECT  1.570 0.870 1.670 4.110 ;
        RECT  1.320 0.870 1.570 1.110 ;
        RECT  1.430 2.920 1.570 4.110 ;
        RECT  1.200 3.710 1.430 4.110 ;
        RECT  0.920 0.730 1.320 1.110 ;
        RECT  1.150 2.240 1.290 2.640 ;
        RECT  0.910 1.390 1.150 3.280 ;
        RECT  0.860 2.880 0.910 3.280 ;
    END
END TLATX1

MACRO TIELO
    CLASS CORE ;
    FOREIGN TIELO 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.270 1.320 1.870 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.490 0.580 5.440 ;
        RECT  0.580 4.640 1.980 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.250 0.400 ;
        RECT  0.250 -0.400 0.490 1.740 ;
        RECT  0.490 -0.400 1.980 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.370 3.210 1.450 3.610 ;
        RECT  1.050 2.980 1.370 3.610 ;
        RECT  0.500 2.980 1.050 3.220 ;
        RECT  0.260 2.170 0.500 3.220 ;
    END
END TIELO

MACRO TIEHI
    CLASS CORE ;
    FOREIGN TIEHI 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 0.880 2.650 ;
        RECT  0.880 2.390 0.900 3.070 ;
        RECT  0.900 2.390 1.120 3.150 ;
        RECT  1.120 2.660 1.210 3.150 ;
        RECT  1.210 2.750 1.300 3.150 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.040 0.580 5.440 ;
        RECT  0.580 4.640 1.980 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.460 0.400 ;
        RECT  0.460 -0.400 0.860 0.560 ;
        RECT  0.860 -0.400 1.980 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  0.610 1.390 1.010 1.790 ;
        RECT  0.500 1.550 0.610 1.790 ;
        RECT  0.260 1.550 0.500 2.390 ;
    END
END TIEHI

MACRO TBUFIXL
    CLASS CORE ;
    FOREIGN TBUFIXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  2.380 3.170 2.720 4.070 ;
        RECT  2.180 1.110 2.720 1.540 ;
        RECT  2.720 1.110 2.960 4.070 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.760 2.150 1.120 2.800 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 2.550 1.520 2.950 ;
        RECT  1.520 2.550 1.780 3.210 ;
        RECT  1.780 2.550 1.800 3.200 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.080 5.440 ;
        RECT  1.080 4.480 1.480 5.440 ;
        RECT  1.480 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.110 0.400 ;
        RECT  1.110 -0.400 1.510 1.310 ;
        RECT  1.510 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.380 2.520 2.440 2.920 ;
        RECT  2.140 1.870 2.380 2.920 ;
        RECT  1.740 1.870 2.140 2.110 ;
        RECT  1.500 1.600 1.740 2.110 ;
        RECT  0.610 1.600 1.500 1.840 ;
        RECT  0.450 3.160 0.780 3.560 ;
        RECT  0.450 0.900 0.610 1.840 ;
        RECT  0.210 0.900 0.450 3.560 ;
    END
END TBUFIXL

MACRO TBUFIX8
    CLASS CORE ;
    FOREIGN TBUFIX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFIXL ;
    SIZE 9.240 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  6.310 2.990 6.710 4.110 ;
        RECT  6.150 1.190 6.710 1.670 ;
        RECT  6.710 2.990 6.810 3.500 ;
        RECT  6.710 1.190 6.810 1.830 ;
        RECT  6.810 1.190 7.850 3.500 ;
        RECT  7.850 1.190 7.970 4.110 ;
        RECT  7.970 1.760 8.250 4.110 ;
        RECT  8.250 1.760 8.370 3.500 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 2.380 2.980 2.660 ;
        RECT  2.980 2.350 3.380 2.750 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.730 1.840 0.860 2.300 ;
        RECT  0.860 1.830 1.110 2.300 ;
        RECT  1.110 1.830 1.120 2.090 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.940 5.440 ;
        RECT  0.940 3.220 1.340 5.440 ;
        RECT  1.340 4.640 2.510 5.440 ;
        RECT  2.510 4.480 2.910 5.440 ;
        RECT  2.910 4.640 5.570 5.440 ;
        RECT  5.570 3.890 5.970 5.440 ;
        RECT  5.970 4.640 7.050 5.440 ;
        RECT  7.050 3.890 7.450 5.440 ;
        RECT  7.450 4.640 8.590 5.440 ;
        RECT  8.590 3.890 8.990 5.440 ;
        RECT  8.990 4.640 9.240 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        RECT  0.940 -0.400 1.340 1.410 ;
        RECT  1.340 -0.400 2.520 0.400 ;
        RECT  2.520 -0.400 2.920 0.560 ;
        RECT  2.920 -0.400 5.510 0.400 ;
        RECT  5.510 -0.400 5.910 0.560 ;
        RECT  5.910 -0.400 6.850 0.400 ;
        RECT  6.850 -0.400 7.250 0.880 ;
        RECT  7.250 -0.400 8.190 0.400 ;
        RECT  8.190 -0.400 8.590 0.880 ;
        RECT  8.590 -0.400 9.240 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.290 2.330 6.530 2.740 ;
        RECT  5.290 2.500 6.290 2.740 ;
        RECT  5.570 0.860 5.810 2.220 ;
        RECT  4.540 0.860 5.570 1.100 ;
        RECT  5.050 1.380 5.290 4.350 ;
        RECT  4.820 1.380 5.050 1.620 ;
        RECT  3.490 4.110 5.050 4.350 ;
        RECT  4.540 2.300 4.570 3.820 ;
        RECT  4.430 0.860 4.540 3.820 ;
        RECT  4.330 0.800 4.430 3.820 ;
        RECT  4.300 0.800 4.330 2.540 ;
        RECT  4.050 3.580 4.330 3.820 ;
        RECT  4.030 0.800 4.300 1.200 ;
        RECT  3.920 2.890 4.040 3.300 ;
        RECT  2.100 0.870 4.030 1.110 ;
        RECT  3.920 1.740 4.020 2.140 ;
        RECT  3.680 1.740 3.920 3.300 ;
        RECT  3.530 1.740 3.680 2.060 ;
        RECT  3.550 3.060 3.680 3.300 ;
        RECT  3.230 3.060 3.550 3.540 ;
        RECT  3.130 1.660 3.530 2.060 ;
        RECT  3.250 3.930 3.490 4.350 ;
        RECT  2.100 3.930 3.250 4.170 ;
        RECT  3.150 3.140 3.230 3.540 ;
        RECT  1.720 0.680 2.100 1.110 ;
        RECT  1.700 3.220 2.100 4.170 ;
        RECT  1.720 1.840 1.800 2.320 ;
        RECT  1.700 0.680 1.720 1.080 ;
        RECT  1.480 1.840 1.720 2.840 ;
        RECT  0.500 2.600 1.480 2.840 ;
        RECT  0.450 1.060 0.580 1.460 ;
        RECT  0.500 3.220 0.580 4.120 ;
        RECT  0.450 2.600 0.500 4.120 ;
        RECT  0.210 1.060 0.450 4.120 ;
        RECT  0.180 1.060 0.210 1.460 ;
        RECT  0.180 3.220 0.210 4.120 ;
    END
END TBUFIX8

MACRO TBUFIX4
    CLASS CORE ;
    FOREIGN TBUFIX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFIXL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  5.270 2.960 5.390 3.940 ;
        RECT  5.390 2.380 5.450 3.940 ;
        RECT  5.450 1.260 5.850 3.940 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.470 2.360 1.480 2.660 ;
        RECT  1.480 2.140 1.880 2.660 ;
        RECT  1.880 2.360 1.890 2.660 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.780 1.840 0.860 2.930 ;
        RECT  0.860 1.830 1.020 2.930 ;
        RECT  1.020 1.830 1.120 2.090 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.010 5.440 ;
        RECT  1.010 4.480 1.410 5.440 ;
        RECT  1.410 4.640 4.510 5.440 ;
        RECT  4.510 3.130 4.910 5.440 ;
        RECT  4.910 4.640 6.040 5.440 ;
        RECT  6.040 4.480 6.440 5.440 ;
        RECT  6.440 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.240 0.400 ;
        RECT  1.240 -0.400 1.640 0.560 ;
        RECT  1.640 -0.400 4.610 0.400 ;
        RECT  4.610 -0.400 5.010 1.360 ;
        RECT  5.010 -0.400 6.040 0.400 ;
        RECT  6.040 -0.400 6.440 0.560 ;
        RECT  6.440 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.920 1.600 5.160 2.020 ;
        RECT  4.170 2.420 5.120 2.660 ;
        RECT  4.310 1.600 4.920 1.840 ;
        RECT  4.070 0.670 4.310 1.840 ;
        RECT  3.790 2.420 4.170 3.800 ;
        RECT  2.980 0.670 4.070 0.910 ;
        RECT  3.770 1.470 3.790 3.800 ;
        RECT  3.550 1.470 3.770 2.660 ;
        RECT  2.620 3.550 3.770 3.790 ;
        RECT  1.930 4.130 3.570 4.370 ;
        RECT  3.260 1.470 3.550 1.870 ;
        RECT  3.030 2.150 3.270 3.270 ;
        RECT  2.980 2.150 3.030 2.390 ;
        RECT  2.740 0.670 2.980 2.390 ;
        RECT  2.460 2.670 2.690 3.070 ;
        RECT  2.210 3.450 2.620 3.790 ;
        RECT  2.220 1.350 2.460 3.170 ;
        RECT  2.060 1.350 2.220 1.790 ;
        RECT  1.790 2.930 2.220 3.170 ;
        RECT  1.480 1.390 2.060 1.790 ;
        RECT  1.690 3.910 1.930 4.370 ;
        RECT  1.380 2.930 1.790 3.260 ;
        RECT  0.960 3.910 1.690 4.150 ;
        RECT  0.720 3.330 0.960 4.150 ;
        RECT  0.500 1.090 0.840 1.490 ;
        RECT  0.560 3.330 0.720 3.730 ;
        RECT  0.500 3.330 0.560 3.570 ;
        RECT  0.260 1.090 0.500 3.570 ;
    END
END TBUFIX4

MACRO TBUFIX3
    CLASS CORE ;
    FOREIGN TBUFIX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFIXL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  5.270 3.030 5.390 4.010 ;
        RECT  5.280 0.690 5.390 1.090 ;
        RECT  5.390 0.690 5.680 4.010 ;
        RECT  5.680 1.820 5.690 4.010 ;
        RECT  5.690 1.820 5.830 2.660 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 2.140 1.520 2.540 ;
        RECT  1.520 2.140 1.780 2.650 ;
        RECT  1.780 2.140 1.880 2.540 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.780 1.840 0.860 2.980 ;
        RECT  0.860 1.830 1.020 2.980 ;
        RECT  1.020 1.830 1.120 2.090 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.980 5.440 ;
        RECT  0.980 4.480 1.380 5.440 ;
        RECT  1.380 4.640 4.510 5.440 ;
        RECT  4.510 2.910 4.910 5.440 ;
        RECT  4.910 4.640 6.030 5.440 ;
        RECT  6.030 3.020 6.430 5.440 ;
        RECT  6.430 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.160 0.400 ;
        RECT  1.160 -0.400 1.560 0.560 ;
        RECT  1.560 -0.400 4.590 0.400 ;
        RECT  4.590 -0.400 4.830 0.940 ;
        RECT  4.830 -0.400 6.030 0.400 ;
        RECT  6.030 -0.400 6.430 1.090 ;
        RECT  6.430 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.720 2.200 5.120 2.600 ;
        RECT  4.710 1.480 5.110 1.880 ;
        RECT  4.150 2.360 4.720 2.600 ;
        RECT  4.290 1.480 4.710 1.720 ;
        RECT  4.050 0.670 4.290 1.720 ;
        RECT  4.150 4.130 4.230 4.370 ;
        RECT  3.990 2.170 4.150 3.340 ;
        RECT  3.830 4.120 4.150 4.370 ;
        RECT  3.030 0.670 4.050 0.910 ;
        RECT  3.910 2.170 3.990 3.790 ;
        RECT  3.760 2.170 3.910 2.410 ;
        RECT  3.750 2.940 3.910 3.790 ;
        RECT  1.930 4.120 3.830 4.360 ;
        RECT  3.520 1.490 3.760 2.410 ;
        RECT  2.620 3.550 3.750 3.790 ;
        RECT  3.310 1.490 3.520 1.890 ;
        RECT  3.220 2.860 3.350 3.280 ;
        RECT  3.030 2.170 3.220 3.280 ;
        RECT  2.980 0.670 3.030 3.280 ;
        RECT  2.790 0.670 2.980 2.410 ;
        RECT  2.510 0.670 2.790 0.930 ;
        RECT  2.430 2.690 2.700 3.090 ;
        RECT  2.210 3.450 2.620 3.790 ;
        RECT  2.430 1.410 2.510 1.810 ;
        RECT  2.190 1.410 2.430 3.170 ;
        RECT  1.480 1.410 2.190 1.810 ;
        RECT  1.790 2.930 2.190 3.170 ;
        RECT  1.690 3.910 1.930 4.360 ;
        RECT  1.380 2.930 1.790 3.260 ;
        RECT  1.000 3.910 1.690 4.150 ;
        RECT  0.760 3.290 1.000 4.150 ;
        RECT  0.500 1.150 0.840 1.550 ;
        RECT  0.600 3.290 0.760 3.690 ;
        RECT  0.500 3.290 0.600 3.530 ;
        RECT  0.440 1.150 0.500 3.530 ;
        RECT  0.260 1.160 0.440 3.530 ;
    END
END TBUFIX3

MACRO TBUFIX2
    CLASS CORE ;
    FOREIGN TBUFIX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFIXL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  2.280 3.560 2.850 3.960 ;
        RECT  2.850 3.560 2.870 3.800 ;
        RECT  2.300 0.970 2.970 1.370 ;
        RECT  2.970 1.130 3.020 1.370 ;
        RECT  2.870 3.430 3.110 3.800 ;
        RECT  3.020 1.130 3.260 2.060 ;
        RECT  3.110 3.430 3.410 3.670 ;
        RECT  3.260 1.820 3.500 2.060 ;
        RECT  3.410 3.220 3.510 3.670 ;
        RECT  3.500 1.820 3.510 2.090 ;
        RECT  3.510 1.820 3.740 3.670 ;
        RECT  3.740 1.830 3.750 3.670 ;
        RECT  3.750 1.830 3.760 2.090 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.770 1.650 0.790 3.100 ;
        RECT  0.790 1.650 1.010 3.210 ;
        RECT  1.010 2.810 1.190 3.210 ;
        RECT  1.010 1.650 2.090 1.890 ;
        RECT  2.090 1.650 2.490 2.050 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.310 2.170 1.470 2.410 ;
        RECT  1.470 2.170 1.710 2.650 ;
        RECT  1.710 2.410 2.810 2.650 ;
        RECT  2.810 2.400 2.840 2.800 ;
        RECT  2.840 2.390 3.100 2.800 ;
        RECT  3.100 2.400 3.210 2.800 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.010 5.440 ;
        RECT  1.010 4.480 1.410 5.440 ;
        RECT  1.410 4.640 3.570 5.440 ;
        RECT  3.570 3.960 3.970 5.440 ;
        RECT  3.970 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.060 0.400 ;
        RECT  1.060 -0.400 1.460 1.370 ;
        RECT  1.460 -0.400 3.540 0.400 ;
        RECT  3.540 -0.400 3.940 1.380 ;
        RECT  3.940 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.040 2.930 2.440 3.260 ;
        RECT  1.730 3.020 2.040 3.260 ;
        RECT  1.490 3.020 1.730 3.780 ;
        RECT  0.570 3.540 1.490 3.780 ;
        RECT  0.490 3.490 0.570 3.890 ;
        RECT  0.250 1.220 0.490 3.890 ;
        RECT  0.160 1.220 0.250 1.640 ;
        RECT  0.170 3.490 0.250 3.890 ;
    END
END TBUFIX2

MACRO TBUFIX20
    CLASS CORE ;
    FOREIGN TBUFIX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFIXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  9.650 2.990 10.090 4.010 ;
        RECT  9.400 1.140 10.720 1.680 ;
        RECT  10.090 2.990 11.230 3.840 ;
        RECT  11.230 2.990 11.630 4.010 ;
        RECT  11.630 2.990 12.090 3.840 ;
        RECT  10.720 1.140 12.090 1.940 ;
        RECT  12.090 1.140 12.770 3.840 ;
        RECT  12.770 1.140 13.170 4.010 ;
        RECT  13.170 1.140 13.650 3.840 ;
        RECT  13.650 2.990 14.310 3.840 ;
        RECT  14.310 2.990 14.710 4.010 ;
        RECT  13.650 1.140 15.340 1.940 ;
        RECT  14.710 2.990 15.850 3.840 ;
        RECT  15.850 2.990 16.250 4.010 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.970 2.390 6.370 2.790 ;
        RECT  6.370 2.550 6.710 2.790 ;
        RECT  6.710 2.550 6.800 3.190 ;
        RECT  6.800 2.550 6.950 3.210 ;
        RECT  6.950 2.950 7.060 3.210 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 1.900 0.860 2.300 ;
        RECT  0.860 1.830 1.120 2.300 ;
        RECT  1.120 1.840 1.280 2.300 ;
        RECT  1.280 1.900 1.640 2.300 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.190 5.440 ;
        RECT  0.190 3.040 0.590 5.440 ;
        RECT  0.590 4.640 1.690 5.440 ;
        RECT  1.690 4.480 2.090 5.440 ;
        RECT  2.090 4.640 3.170 5.440 ;
        RECT  3.170 4.120 3.570 5.440 ;
        RECT  3.570 4.640 4.660 5.440 ;
        RECT  4.660 4.480 5.060 5.440 ;
        RECT  5.060 4.640 8.950 5.440 ;
        RECT  8.950 4.250 9.350 5.440 ;
        RECT  9.350 4.640 10.430 5.440 ;
        RECT  10.430 4.120 10.830 5.440 ;
        RECT  10.830 4.640 11.970 5.440 ;
        RECT  11.970 4.120 12.370 5.440 ;
        RECT  12.370 4.640 13.510 5.440 ;
        RECT  13.510 4.120 13.910 5.440 ;
        RECT  13.910 4.640 15.050 5.440 ;
        RECT  15.050 4.120 15.450 5.440 ;
        RECT  15.450 4.640 16.590 5.440 ;
        RECT  16.590 4.090 16.990 5.440 ;
        RECT  16.990 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.370 0.400 ;
        RECT  0.370 -0.400 0.770 1.530 ;
        RECT  0.770 -0.400 1.980 0.400 ;
        RECT  1.980 -0.400 2.380 0.560 ;
        RECT  2.380 -0.400 3.380 0.400 ;
        RECT  3.380 -0.400 3.780 1.040 ;
        RECT  3.780 -0.400 4.720 0.400 ;
        RECT  4.720 -0.400 5.120 0.560 ;
        RECT  5.120 -0.400 8.760 0.400 ;
        RECT  8.760 -0.400 9.160 0.560 ;
        RECT  9.160 -0.400 10.130 0.400 ;
        RECT  10.130 -0.400 10.530 0.870 ;
        RECT  10.530 -0.400 11.470 0.400 ;
        RECT  11.470 -0.400 11.870 0.870 ;
        RECT  11.870 -0.400 12.810 0.400 ;
        RECT  12.810 -0.400 13.210 0.870 ;
        RECT  13.210 -0.400 14.160 0.400 ;
        RECT  14.160 -0.400 14.560 0.870 ;
        RECT  14.560 -0.400 15.540 0.400 ;
        RECT  15.540 -0.400 15.940 0.870 ;
        RECT  15.940 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.560 2.320 11.610 2.730 ;
        RECT  9.390 2.480 10.560 2.720 ;
        RECT  8.910 1.950 10.200 2.190 ;
        RECT  9.150 2.480 9.390 4.010 ;
        RECT  8.430 3.770 9.150 4.010 ;
        RECT  8.670 0.860 8.910 3.430 ;
        RECT  7.470 0.860 8.670 1.100 ;
        RECT  7.680 3.190 8.670 3.430 ;
        RECT  8.190 3.770 8.430 4.350 ;
        RECT  8.180 1.390 8.340 1.630 ;
        RECT  8.030 3.820 8.190 4.350 ;
        RECT  7.940 1.390 8.180 2.150 ;
        RECT  5.020 3.820 8.030 4.060 ;
        RECT  7.910 1.910 7.940 2.150 ;
        RECT  7.510 1.910 7.910 2.700 ;
        RECT  7.440 3.110 7.680 3.510 ;
        RECT  5.610 1.910 7.510 2.150 ;
        RECT  7.060 0.670 7.470 1.100 ;
        RECT  5.940 0.670 7.060 0.910 ;
        RECT  6.300 1.220 6.700 1.620 ;
        RECT  5.020 1.380 6.300 1.620 ;
        RECT  5.620 0.670 5.940 1.100 ;
        RECT  5.610 3.100 5.880 3.500 ;
        RECT  4.450 0.860 5.620 1.100 ;
        RECT  5.480 1.910 5.610 3.500 ;
        RECT  5.370 1.910 5.480 3.420 ;
        RECT  4.780 1.380 5.020 4.060 ;
        RECT  2.430 3.320 4.780 3.720 ;
        RECT  4.210 0.860 4.450 1.720 ;
        RECT  3.180 2.010 4.440 2.410 ;
        RECT  2.710 1.320 4.210 1.720 ;
        RECT  2.370 2.000 3.180 2.410 ;
        RECT  2.130 1.310 2.370 2.900 ;
        RECT  1.580 1.310 2.130 1.550 ;
        RECT  1.310 2.660 2.130 2.900 ;
        RECT  1.180 1.150 1.580 1.550 ;
        RECT  0.910 2.660 1.310 3.860 ;
    END
END TBUFIX20

MACRO TBUFIX1
    CLASS CORE ;
    FOREIGN TBUFIX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFIXL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  2.420 3.260 2.750 4.160 ;
        RECT  2.750 3.220 2.800 4.160 ;
        RECT  2.180 1.030 2.800 1.540 ;
        RECT  2.800 1.030 2.820 4.160 ;
        RECT  2.820 1.030 3.040 3.520 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.730 1.850 1.140 2.110 ;
        RECT  1.140 1.850 1.520 2.090 ;
        RECT  1.520 1.820 2.480 2.100 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 1.120 2.650 ;
        RECT  1.120 2.410 1.210 2.650 ;
        RECT  1.210 2.410 1.450 2.890 ;
        RECT  1.450 2.490 1.530 2.890 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.070 5.440 ;
        RECT  1.070 4.480 1.470 5.440 ;
        RECT  1.470 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.040 0.400 ;
        RECT  1.040 -0.400 1.110 0.560 ;
        RECT  1.110 -0.400 1.510 1.440 ;
        RECT  1.510 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.090 2.570 2.490 2.970 ;
        RECT  2.050 2.730 2.090 2.970 ;
        RECT  1.810 2.730 2.050 3.420 ;
        RECT  0.590 3.180 1.810 3.420 ;
        RECT  0.450 1.180 0.590 1.580 ;
        RECT  0.450 3.180 0.590 3.610 ;
        RECT  0.210 1.180 0.450 3.610 ;
        RECT  0.190 1.180 0.210 1.580 ;
        RECT  0.190 3.210 0.210 3.610 ;
    END
END TBUFIX1

MACRO TBUFIX16
    CLASS CORE ;
    FOREIGN TBUFIX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFIXL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  9.110 2.990 9.550 4.190 ;
        RECT  8.910 1.140 10.160 1.680 ;
        RECT  9.550 2.990 10.670 3.840 ;
        RECT  10.670 2.990 10.690 4.060 ;
        RECT  10.690 2.990 11.090 4.190 ;
        RECT  11.090 2.990 11.110 4.060 ;
        RECT  11.110 2.990 11.430 3.840 ;
        RECT  10.160 1.140 11.430 1.940 ;
        RECT  11.430 1.140 12.230 3.840 ;
        RECT  12.230 1.140 12.630 4.190 ;
        RECT  12.630 1.140 12.990 3.840 ;
        RECT  12.990 1.140 13.510 1.940 ;
        RECT  12.990 2.990 13.770 3.840 ;
        RECT  13.770 2.990 14.170 4.190 ;
        RECT  14.170 2.990 14.210 3.840 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.620 1.940 5.780 2.340 ;
        RECT  5.780 1.860 6.020 2.340 ;
        RECT  6.020 1.860 6.140 2.100 ;
        RECT  6.140 1.830 6.390 2.100 ;
        RECT  6.390 1.830 6.400 2.090 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.960 1.900 1.520 2.300 ;
        RECT  1.520 1.830 1.780 2.300 ;
        RECT  1.780 1.900 1.920 2.300 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.290 5.440 ;
        RECT  0.290 2.800 0.690 5.440 ;
        RECT  0.690 4.640 1.810 5.440 ;
        RECT  1.810 4.480 2.210 5.440 ;
        RECT  2.210 4.640 3.280 5.440 ;
        RECT  3.280 4.120 3.680 5.440 ;
        RECT  3.680 4.640 4.930 5.440 ;
        RECT  4.930 4.080 5.610 5.440 ;
        RECT  5.610 4.640 8.370 5.440 ;
        RECT  8.370 4.060 8.770 5.440 ;
        RECT  8.770 4.640 9.870 5.440 ;
        RECT  9.870 4.160 10.270 5.440 ;
        RECT  10.270 4.640 11.430 5.440 ;
        RECT  11.430 4.110 11.830 5.440 ;
        RECT  11.830 4.640 12.970 5.440 ;
        RECT  12.970 4.110 13.370 5.440 ;
        RECT  13.370 4.640 14.490 5.440 ;
        RECT  14.490 4.110 14.890 5.440 ;
        RECT  14.890 4.640 15.180 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.790 0.400 ;
        RECT  0.790 -0.400 1.190 1.440 ;
        RECT  1.190 -0.400 2.240 0.400 ;
        RECT  2.240 -0.400 2.640 0.560 ;
        RECT  2.640 -0.400 3.590 0.400 ;
        RECT  3.590 -0.400 3.990 0.900 ;
        RECT  3.990 -0.400 6.640 0.400 ;
        RECT  6.640 -0.400 7.040 0.560 ;
        RECT  7.040 -0.400 8.310 0.400 ;
        RECT  8.310 -0.400 8.710 0.560 ;
        RECT  8.710 -0.400 9.650 0.400 ;
        RECT  9.650 -0.400 10.050 0.870 ;
        RECT  10.050 -0.400 10.990 0.400 ;
        RECT  10.990 -0.400 11.390 0.870 ;
        RECT  11.390 -0.400 12.330 0.400 ;
        RECT  12.330 -0.400 12.730 0.870 ;
        RECT  12.730 -0.400 13.700 0.400 ;
        RECT  13.700 -0.400 14.100 0.870 ;
        RECT  14.100 -0.400 15.180 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.560 2.410 10.980 2.730 ;
        RECT  10.000 2.410 10.560 2.720 ;
        RECT  8.710 2.480 10.000 2.720 ;
        RECT  8.550 1.950 9.710 2.190 ;
        RECT  8.470 2.480 8.710 3.540 ;
        RECT  8.310 0.860 8.550 2.190 ;
        RECT  8.080 3.300 8.470 3.540 ;
        RECT  6.200 0.860 8.310 1.100 ;
        RECT  8.130 1.950 8.310 2.190 ;
        RECT  7.890 1.950 8.130 3.010 ;
        RECT  7.840 3.300 8.080 4.350 ;
        RECT  7.550 1.380 7.960 1.670 ;
        RECT  7.520 2.770 7.890 3.010 ;
        RECT  6.260 4.110 7.840 4.350 ;
        RECT  7.380 1.430 7.550 1.670 ;
        RECT  7.280 2.770 7.520 3.510 ;
        RECT  7.060 1.430 7.380 1.890 ;
        RECT  7.200 3.270 7.280 3.510 ;
        RECT  6.800 3.270 7.200 3.670 ;
        RECT  7.000 1.490 7.060 1.890 ;
        RECT  6.980 1.490 7.000 2.890 ;
        RECT  6.760 1.650 6.980 2.890 ;
        RECT  6.530 2.650 6.760 2.890 ;
        RECT  6.130 2.650 6.530 3.110 ;
        RECT  6.020 3.550 6.260 4.350 ;
        RECT  6.040 0.860 6.200 1.370 ;
        RECT  5.390 2.870 6.130 3.110 ;
        RECT  5.800 0.670 6.040 1.370 ;
        RECT  4.410 3.550 6.020 3.790 ;
        RECT  4.670 0.670 5.800 0.910 ;
        RECT  5.280 1.190 5.440 1.520 ;
        RECT  4.990 2.870 5.390 3.270 ;
        RECT  5.040 1.190 5.280 2.570 ;
        RECT  4.410 2.330 5.040 2.570 ;
        RECT  4.590 0.670 4.670 1.610 ;
        RECT  4.430 0.670 4.590 1.640 ;
        RECT  4.270 1.210 4.430 1.640 ;
        RECT  4.170 2.330 4.410 3.790 ;
        RECT  2.980 1.400 4.270 1.640 ;
        RECT  4.070 3.180 4.170 3.790 ;
        RECT  2.530 3.180 4.070 3.580 ;
        RECT  2.410 1.920 3.660 2.320 ;
        RECT  2.170 1.310 2.410 2.900 ;
        RECT  1.950 1.310 2.170 1.550 ;
        RECT  1.410 2.660 2.170 2.900 ;
        RECT  1.550 1.150 1.950 1.550 ;
        RECT  1.010 2.660 1.410 3.760 ;
    END
END TBUFIX16

MACRO TBUFIX12
    CLASS CORE ;
    FOREIGN TBUFIX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFIXL ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  8.190 1.140 9.460 1.680 ;
        RECT  8.130 2.990 9.710 3.670 ;
        RECT  9.710 2.990 10.110 4.000 ;
        RECT  9.460 1.140 10.110 1.820 ;
        RECT  10.110 1.140 11.170 3.670 ;
        RECT  11.170 1.140 11.530 4.000 ;
        RECT  11.530 1.200 11.650 4.000 ;
        RECT  11.650 1.200 11.670 3.630 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 1.830 4.270 2.090 ;
        RECT  4.270 1.830 4.420 2.490 ;
        RECT  4.420 1.850 4.510 2.490 ;
        RECT  4.510 2.250 4.940 2.490 ;
        RECT  4.940 2.250 5.340 2.650 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.390 1.840 1.520 2.300 ;
        RECT  1.520 1.830 1.770 2.300 ;
        RECT  1.770 1.830 1.780 2.090 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.410 5.440 ;
        RECT  1.410 4.180 1.810 5.440 ;
        RECT  1.810 4.640 2.730 5.440 ;
        RECT  2.730 4.170 3.130 5.440 ;
        RECT  3.130 4.640 4.130 5.440 ;
        RECT  4.130 4.080 4.790 5.440 ;
        RECT  4.790 4.640 7.430 5.440 ;
        RECT  7.430 4.140 7.830 5.440 ;
        RECT  7.830 4.640 8.910 5.440 ;
        RECT  8.910 3.940 9.310 5.440 ;
        RECT  9.310 4.640 10.450 5.440 ;
        RECT  10.450 3.940 10.850 5.440 ;
        RECT  10.850 4.640 11.970 5.440 ;
        RECT  11.970 3.940 12.370 5.440 ;
        RECT  12.370 4.640 12.540 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.600 0.400 ;
        RECT  1.600 -0.400 2.000 1.570 ;
        RECT  2.000 -0.400 3.160 0.400 ;
        RECT  3.160 -0.400 3.560 1.010 ;
        RECT  3.560 -0.400 5.390 0.400 ;
        RECT  5.390 -0.400 5.790 0.560 ;
        RECT  5.790 -0.400 7.590 0.400 ;
        RECT  7.590 -0.400 7.990 0.560 ;
        RECT  7.990 -0.400 8.930 0.400 ;
        RECT  8.930 -0.400 9.330 0.870 ;
        RECT  9.330 -0.400 10.270 0.400 ;
        RECT  10.270 -0.400 10.670 0.870 ;
        RECT  10.670 -0.400 11.610 0.400 ;
        RECT  11.610 -0.400 12.010 0.870 ;
        RECT  12.010 -0.400 12.540 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  9.570 2.390 9.650 2.630 ;
        RECT  9.220 2.390 9.570 2.720 ;
        RECT  7.370 2.480 9.220 2.720 ;
        RECT  7.910 1.940 8.530 2.180 ;
        RECT  7.670 0.860 7.910 2.180 ;
        RECT  6.660 0.860 7.670 1.100 ;
        RECT  7.130 1.380 7.370 2.720 ;
        RECT  6.900 1.380 7.130 1.620 ;
        RECT  7.060 2.480 7.130 2.720 ;
        RECT  6.820 2.480 7.060 4.350 ;
        RECT  5.390 4.110 6.820 4.350 ;
        RECT  6.580 0.670 6.660 1.100 ;
        RECT  6.340 0.670 6.580 3.830 ;
        RECT  6.260 0.670 6.340 1.110 ;
        RECT  5.870 3.590 6.340 3.830 ;
        RECT  4.360 0.870 6.260 1.110 ;
        RECT  5.940 1.730 6.100 2.140 ;
        RECT  5.700 1.730 5.940 3.300 ;
        RECT  5.330 1.730 5.700 1.970 ;
        RECT  4.590 3.030 5.700 3.270 ;
        RECT  5.150 3.550 5.390 4.350 ;
        RECT  4.930 1.510 5.330 1.970 ;
        RECT  3.740 3.550 5.150 3.790 ;
        RECT  4.190 2.870 4.590 3.270 ;
        RECT  3.960 0.680 4.360 1.580 ;
        RECT  2.760 1.340 3.960 1.580 ;
        RECT  3.340 3.320 3.740 3.790 ;
        RECT  2.020 3.320 3.340 3.720 ;
        RECT  2.370 1.920 3.110 2.320 ;
        RECT  2.440 0.670 2.760 1.580 ;
        RECT  2.360 0.670 2.440 1.570 ;
        RECT  2.130 1.920 2.370 2.840 ;
        RECT  0.930 2.600 2.130 2.840 ;
        RECT  0.840 0.640 1.240 1.540 ;
        RECT  0.800 2.600 0.930 4.400 ;
        RECT  0.800 1.300 0.840 1.540 ;
        RECT  0.560 1.300 0.800 4.400 ;
        RECT  0.530 2.900 0.560 4.400 ;
    END
END TBUFIX12

MACRO TBUFXL
    CLASS CORE ;
    FOREIGN TBUFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  4.250 3.170 4.720 3.570 ;
        RECT  4.360 1.190 4.720 1.590 ;
        RECT  4.720 1.190 5.120 3.570 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.800 1.760 1.360 2.160 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.180 2.450 3.410 2.850 ;
        RECT  3.410 2.450 3.500 3.190 ;
        RECT  3.500 2.450 3.580 3.210 ;
        RECT  3.580 2.610 3.650 3.210 ;
        RECT  3.650 2.950 3.760 3.210 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.090 5.440 ;
        RECT  1.090 4.480 1.490 5.440 ;
        RECT  1.490 4.640 3.400 5.440 ;
        RECT  3.400 4.480 3.800 5.440 ;
        RECT  3.800 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.120 0.400 ;
        RECT  1.120 -0.400 1.520 0.560 ;
        RECT  1.520 -0.400 3.960 0.400 ;
        RECT  3.960 -0.400 4.360 0.560 ;
        RECT  4.360 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.450 4.010 4.460 4.250 ;
        RECT  4.060 3.940 4.450 4.250 ;
        RECT  4.040 1.860 4.440 2.260 ;
        RECT  3.060 3.940 4.060 4.180 ;
        RECT  3.680 1.860 4.040 2.100 ;
        RECT  3.440 0.680 3.680 2.100 ;
        RECT  2.140 0.680 3.440 0.920 ;
        RECT  2.890 1.390 3.100 1.790 ;
        RECT  2.890 3.170 3.060 4.180 ;
        RECT  2.650 1.390 2.890 4.180 ;
        RECT  0.600 3.940 2.650 4.180 ;
        RECT  1.900 0.680 2.140 3.570 ;
        RECT  1.740 3.170 1.900 3.570 ;
        RECT  1.320 1.020 1.560 1.420 ;
        RECT  1.320 2.480 1.560 2.880 ;
        RECT  0.620 1.100 1.320 1.340 ;
        RECT  0.610 2.560 1.320 2.800 ;
        RECT  0.420 0.670 0.620 1.340 ;
        RECT  0.420 2.560 0.610 3.510 ;
        RECT  0.200 3.890 0.600 4.290 ;
        RECT  0.180 0.670 0.420 3.510 ;
    END
END TBUFXL

MACRO TBUFX8
    CLASS CORE ;
    FOREIGN TBUFX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFXL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  4.730 3.010 5.130 4.070 ;
        RECT  5.130 3.010 5.610 3.690 ;
        RECT  5.610 2.940 6.000 3.690 ;
        RECT  6.000 1.140 6.250 3.690 ;
        RECT  6.250 1.140 6.650 4.070 ;
        RECT  6.650 1.140 7.720 3.690 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.730 2.110 1.160 2.650 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 2.680 1.720 3.450 ;
        RECT  1.720 3.080 1.870 3.450 ;
        RECT  1.870 3.210 2.940 3.450 ;
        RECT  2.940 2.420 3.180 3.450 ;
        RECT  3.180 2.420 3.280 2.660 ;
        RECT  3.280 2.190 3.520 2.660 ;
        RECT  3.520 2.190 3.680 2.650 ;
        RECT  3.680 2.390 3.760 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.940 5.440 ;
        RECT  0.940 4.260 1.340 5.440 ;
        RECT  1.340 4.640 3.910 5.440 ;
        RECT  3.910 4.250 4.310 5.440 ;
        RECT  4.310 4.640 5.490 5.440 ;
        RECT  5.490 3.960 5.890 5.440 ;
        RECT  5.890 4.640 7.010 5.440 ;
        RECT  7.010 3.960 7.410 5.440 ;
        RECT  7.410 4.640 8.580 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.050 0.400 ;
        RECT  1.050 -0.400 1.450 1.310 ;
        RECT  1.450 -0.400 3.530 0.400 ;
        RECT  3.530 -0.400 3.770 0.870 ;
        RECT  3.770 -0.400 5.090 0.400 ;
        RECT  5.090 -0.400 5.490 1.370 ;
        RECT  5.490 -0.400 6.620 0.400 ;
        RECT  6.620 -0.400 7.020 0.800 ;
        RECT  7.020 -0.400 8.000 0.400 ;
        RECT  8.000 -0.400 8.400 0.800 ;
        RECT  8.400 -0.400 8.580 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.480 1.640 5.720 2.120 ;
        RECT  4.840 1.640 5.480 1.880 ;
        RECT  4.360 2.150 4.880 2.550 ;
        RECT  4.600 1.150 4.840 1.880 ;
        RECT  4.570 1.150 4.600 1.390 ;
        RECT  4.170 1.050 4.570 1.390 ;
        RECT  4.120 1.670 4.360 3.970 ;
        RECT  3.290 1.150 4.170 1.390 ;
        RECT  2.810 1.670 4.120 1.910 ;
        RECT  3.530 3.730 4.120 3.970 ;
        RECT  3.290 3.730 3.530 4.160 ;
        RECT  3.050 0.670 3.290 1.390 ;
        RECT  2.160 3.920 3.290 4.160 ;
        RECT  2.170 0.670 3.050 0.910 ;
        RECT  2.570 1.200 2.810 1.910 ;
        RECT  2.440 2.690 2.660 2.930 ;
        RECT  2.200 2.190 2.440 2.930 ;
        RECT  2.170 2.190 2.200 2.430 ;
        RECT  1.930 0.670 2.170 2.430 ;
        RECT  1.990 3.920 2.160 4.300 ;
        RECT  1.750 3.730 1.990 4.300 ;
        RECT  1.770 1.070 1.930 1.310 ;
        RECT  0.570 3.730 1.750 3.970 ;
        RECT  1.440 1.590 1.680 2.210 ;
        RECT  0.410 1.590 1.440 1.830 ;
        RECT  0.410 0.870 0.570 1.270 ;
        RECT  0.170 3.720 0.570 4.120 ;
        RECT  0.410 2.790 0.490 3.190 ;
        RECT  0.170 0.870 0.410 3.190 ;
    END
END TBUFX8

MACRO TBUFX4
    CLASS CORE ;
    FOREIGN TBUFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFXL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  4.570 0.920 4.730 1.320 ;
        RECT  4.610 3.460 4.770 4.360 ;
        RECT  4.730 0.920 4.770 2.660 ;
        RECT  4.770 0.920 5.050 4.360 ;
        RECT  5.050 1.260 5.090 4.360 ;
        RECT  5.090 1.260 5.170 2.660 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 3.510 0.210 3.770 ;
        RECT  0.210 2.990 0.490 3.770 ;
        RECT  0.490 3.080 0.500 3.770 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 2.130 3.690 2.530 ;
        RECT  3.690 2.130 3.740 3.180 ;
        RECT  3.740 2.290 3.930 3.180 ;
        RECT  3.930 2.940 4.160 3.180 ;
        RECT  4.160 2.940 4.400 3.210 ;
        RECT  4.400 2.950 4.420 3.210 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.340 5.440 ;
        RECT  1.340 4.480 1.740 5.440 ;
        RECT  1.740 4.640 3.850 5.440 ;
        RECT  3.850 3.520 4.250 5.440 ;
        RECT  4.250 4.640 5.370 5.440 ;
        RECT  5.370 3.180 5.770 5.440 ;
        RECT  5.770 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.460 0.400 ;
        RECT  0.460 -0.400 0.860 0.560 ;
        RECT  0.860 -0.400 3.810 0.400 ;
        RECT  3.810 -0.400 4.210 1.320 ;
        RECT  4.210 -0.400 5.330 0.400 ;
        RECT  5.330 -0.400 5.730 0.940 ;
        RECT  5.730 -0.400 5.940 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.220 1.610 4.460 2.630 ;
        RECT  3.150 1.610 4.220 1.850 ;
        RECT  3.290 1.080 3.450 1.320 ;
        RECT  3.170 2.820 3.410 4.180 ;
        RECT  3.050 0.670 3.290 1.320 ;
        RECT  3.150 2.820 3.170 3.060 ;
        RECT  1.910 3.940 3.170 4.180 ;
        RECT  2.910 1.610 3.150 3.060 ;
        RECT  2.480 0.670 3.050 0.920 ;
        RECT  2.200 1.610 2.910 1.850 ;
        RECT  2.630 3.420 2.730 3.660 ;
        RECT  2.390 2.150 2.630 3.660 ;
        RECT  2.210 0.680 2.480 0.920 ;
        RECT  1.920 2.150 2.390 2.390 ;
        RECT  2.330 3.420 2.390 3.660 ;
        RECT  1.970 0.680 2.210 1.310 ;
        RECT  1.060 2.690 2.110 3.090 ;
        RECT  1.920 1.070 1.970 1.310 ;
        RECT  1.680 1.070 1.920 2.390 ;
        RECT  1.670 3.510 1.910 4.180 ;
        RECT  1.160 1.410 1.400 1.820 ;
        RECT  1.060 1.420 1.160 1.820 ;
        RECT  0.840 1.420 1.060 4.290 ;
        RECT  0.820 1.280 0.840 4.290 ;
        RECT  0.440 1.280 0.820 1.680 ;
        RECT  0.170 4.050 0.820 4.290 ;
    END
END TBUFX4

MACRO TBUFX3
    CLASS CORE ;
    FOREIGN TBUFX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFXL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  4.090 3.160 4.290 3.600 ;
        RECT  4.290 2.940 4.730 3.600 ;
        RECT  4.320 1.120 4.730 1.560 ;
        RECT  4.730 1.120 5.170 3.600 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.730 1.830 1.150 2.300 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.090 2.420 3.330 2.860 ;
        RECT  3.330 2.420 3.500 2.660 ;
        RECT  3.500 2.390 3.740 2.660 ;
        RECT  3.740 2.390 3.760 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.060 5.440 ;
        RECT  1.060 4.480 1.460 5.440 ;
        RECT  1.460 4.640 3.440 5.440 ;
        RECT  3.440 4.480 3.840 5.440 ;
        RECT  3.840 4.640 4.840 5.440 ;
        RECT  4.840 4.480 5.240 5.440 ;
        RECT  5.240 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.060 0.400 ;
        RECT  1.060 -0.400 1.460 0.560 ;
        RECT  1.460 -0.400 3.600 0.400 ;
        RECT  3.600 -0.400 3.610 0.670 ;
        RECT  3.610 -0.400 4.010 0.870 ;
        RECT  4.010 -0.400 4.020 0.670 ;
        RECT  4.020 -0.400 5.070 0.400 ;
        RECT  5.070 -0.400 5.470 0.560 ;
        RECT  5.470 -0.400 5.940 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.440 2.430 5.680 4.180 ;
        RECT  2.870 3.940 5.440 4.180 ;
        RECT  3.330 1.830 4.440 2.070 ;
        RECT  3.090 0.730 3.330 2.070 ;
        RECT  2.280 0.730 3.090 0.970 ;
        RECT  2.800 3.780 2.870 4.180 ;
        RECT  2.800 1.620 2.810 2.020 ;
        RECT  2.560 1.620 2.800 4.180 ;
        RECT  2.470 3.780 2.560 4.180 ;
        RECT  0.580 3.940 2.470 4.180 ;
        RECT  2.040 0.730 2.280 3.500 ;
        RECT  1.650 3.260 2.040 3.500 ;
        RECT  1.520 1.110 1.760 1.530 ;
        RECT  1.520 2.580 1.760 2.980 ;
        RECT  0.580 1.290 1.520 1.530 ;
        RECT  0.580 2.740 1.520 2.980 ;
        RECT  0.410 0.940 0.580 1.530 ;
        RECT  0.410 2.740 0.580 3.460 ;
        RECT  0.180 3.940 0.580 4.360 ;
        RECT  0.170 0.940 0.410 3.460 ;
    END
END TBUFX3

MACRO TBUFX2
    CLASS CORE ;
    FOREIGN TBUFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFXL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  4.340 3.130 4.620 3.530 ;
        RECT  4.380 1.230 4.620 1.630 ;
        RECT  4.620 1.230 4.780 3.530 ;
        RECT  4.780 1.310 4.860 3.530 ;
        RECT  4.860 1.830 5.080 2.090 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 0.870 2.090 ;
        RECT  0.870 1.830 1.120 2.290 ;
        RECT  1.120 1.890 1.300 2.290 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.050 2.400 3.410 2.800 ;
        RECT  3.410 2.400 3.450 3.190 ;
        RECT  3.450 2.560 3.500 3.190 ;
        RECT  3.500 2.560 3.650 3.210 ;
        RECT  3.650 2.950 3.760 3.210 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.120 5.440 ;
        RECT  1.120 4.480 1.520 5.440 ;
        RECT  1.520 4.640 3.490 5.440 ;
        RECT  3.490 4.480 3.890 5.440 ;
        RECT  3.890 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.120 0.400 ;
        RECT  1.120 -0.400 1.520 0.560 ;
        RECT  1.520 -0.400 3.540 0.400 ;
        RECT  3.540 -0.400 3.940 0.560 ;
        RECT  3.940 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.510 4.130 5.060 4.370 ;
        RECT  4.240 3.870 4.510 4.370 ;
        RECT  2.990 3.870 4.240 4.110 ;
        RECT  3.900 1.720 4.060 2.120 ;
        RECT  3.660 0.860 3.900 2.120 ;
        RECT  3.100 0.860 3.660 1.100 ;
        RECT  2.080 0.690 3.100 1.100 ;
        RECT  2.650 3.210 2.990 4.110 ;
        RECT  2.650 1.510 2.830 1.910 ;
        RECT  2.410 1.510 2.650 4.110 ;
        RECT  0.600 3.870 2.410 4.110 ;
        RECT  2.030 0.690 2.080 3.540 ;
        RECT  1.840 0.860 2.030 3.540 ;
        RECT  1.670 3.300 1.840 3.540 ;
        RECT  1.320 1.150 1.560 1.550 ;
        RECT  1.320 2.610 1.560 3.010 ;
        RECT  0.600 1.230 1.320 1.470 ;
        RECT  0.600 2.690 1.320 2.930 ;
        RECT  0.430 0.780 0.600 1.470 ;
        RECT  0.430 2.690 0.600 3.470 ;
        RECT  0.200 3.870 0.600 4.350 ;
        RECT  0.190 0.780 0.430 3.470 ;
    END
END TBUFX2

MACRO TBUFX20
    CLASS CORE ;
    FOREIGN TBUFX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  9.110 2.660 10.670 3.460 ;
        RECT  10.670 2.660 10.770 3.640 ;
        RECT  9.660 1.140 10.770 1.940 ;
        RECT  10.770 1.140 12.330 3.840 ;
        RECT  12.330 2.660 12.430 3.640 ;
        RECT  12.330 1.140 15.380 1.940 ;
        RECT  15.380 1.140 15.390 1.540 ;
        RECT  12.430 2.660 15.750 3.460 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.950 0.210 3.210 ;
        RECT  0.210 2.260 0.450 3.210 ;
        RECT  0.450 2.950 0.460 3.210 ;
        RECT  0.450 2.260 0.790 2.500 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.560 1.840 6.800 2.240 ;
        RECT  6.800 1.830 7.060 2.240 ;
        RECT  7.060 1.840 7.660 2.240 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 3.690 5.440 ;
        RECT  3.690 4.480 4.090 5.440 ;
        RECT  4.090 4.640 5.130 5.440 ;
        RECT  5.130 3.720 5.530 5.440 ;
        RECT  5.530 4.640 6.710 5.440 ;
        RECT  6.710 3.960 7.110 5.440 ;
        RECT  7.110 4.640 8.340 5.440 ;
        RECT  8.340 3.470 8.740 5.440 ;
        RECT  8.740 4.640 9.940 5.440 ;
        RECT  9.940 3.910 10.340 5.440 ;
        RECT  10.340 4.640 11.460 5.440 ;
        RECT  11.460 4.280 11.860 5.440 ;
        RECT  11.860 4.640 13.030 5.440 ;
        RECT  13.030 3.900 13.430 5.440 ;
        RECT  13.430 4.640 14.560 5.440 ;
        RECT  14.560 3.900 14.960 5.440 ;
        RECT  14.960 4.640 15.930 5.440 ;
        RECT  15.930 3.900 16.330 5.440 ;
        RECT  16.330 4.640 16.500 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.930 0.400 ;
        RECT  0.930 -0.400 1.330 1.460 ;
        RECT  1.330 -0.400 2.430 0.400 ;
        RECT  2.430 -0.400 2.830 1.330 ;
        RECT  2.830 -0.400 5.400 0.400 ;
        RECT  5.400 -0.400 5.800 0.870 ;
        RECT  5.800 -0.400 6.680 0.400 ;
        RECT  6.680 -0.400 7.080 0.870 ;
        RECT  7.080 -0.400 10.280 0.400 ;
        RECT  10.280 -0.400 10.680 0.870 ;
        RECT  10.680 -0.400 11.620 0.400 ;
        RECT  11.620 -0.400 12.020 0.870 ;
        RECT  12.020 -0.400 12.960 0.400 ;
        RECT  12.960 -0.400 13.360 0.870 ;
        RECT  13.360 -0.400 14.300 0.400 ;
        RECT  14.300 -0.400 14.700 0.870 ;
        RECT  14.700 -0.400 15.620 0.400 ;
        RECT  15.620 -0.400 16.020 0.870 ;
        RECT  16.020 -0.400 16.500 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  8.970 1.150 9.370 1.800 ;
        RECT  7.770 1.150 8.970 1.550 ;
        RECT  8.300 2.070 8.800 3.210 ;
        RECT  4.720 2.710 8.300 3.210 ;
        RECT  5.130 1.140 7.770 1.560 ;
        RECT  5.120 0.670 5.130 1.560 ;
        RECT  4.720 0.670 5.120 1.630 ;
        RECT  4.710 0.670 4.720 1.560 ;
        RECT  4.350 2.710 4.720 3.840 ;
        RECT  3.600 0.670 4.710 1.090 ;
        RECT  3.950 1.390 4.350 3.840 ;
        RECT  2.750 3.420 3.950 3.840 ;
        RECT  3.590 0.670 3.600 1.220 ;
        RECT  3.350 0.670 3.590 2.020 ;
        RECT  3.190 0.670 3.350 3.150 ;
        RECT  3.180 0.670 3.190 1.220 ;
        RECT  2.950 1.610 3.190 3.150 ;
        RECT  2.070 1.610 2.950 1.950 ;
        RECT  1.710 2.750 2.950 3.150 ;
        RECT  2.740 3.420 2.750 3.880 ;
        RECT  2.340 3.420 2.740 4.080 ;
        RECT  1.370 2.230 2.550 2.470 ;
        RECT  2.330 3.420 2.340 3.880 ;
        RECT  1.670 1.330 2.070 1.950 ;
        RECT  1.660 1.360 1.670 1.950 ;
        RECT  1.130 1.740 1.370 3.900 ;
        RECT  0.570 1.740 1.130 1.980 ;
        RECT  0.970 3.000 1.130 3.900 ;
        RECT  0.170 1.320 0.570 1.980 ;
    END
END TBUFX20

MACRO TBUFX1
    CLASS CORE ;
    FOREIGN TBUFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFXL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  4.260 3.130 4.480 3.530 ;
        RECT  4.260 1.140 4.480 1.540 ;
        RECT  4.480 1.140 4.660 3.530 ;
        RECT  4.660 1.170 4.720 3.530 ;
        RECT  4.720 1.820 5.080 3.220 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.780 1.830 1.180 2.290 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.980 2.400 3.380 2.800 ;
        RECT  3.380 2.560 3.410 2.800 ;
        RECT  3.410 2.560 3.500 3.190 ;
        RECT  3.500 2.560 3.650 3.210 ;
        RECT  3.650 2.950 3.760 3.210 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.120 5.440 ;
        RECT  1.120 4.480 1.520 5.440 ;
        RECT  1.520 4.640 3.430 5.440 ;
        RECT  3.430 4.480 3.830 5.440 ;
        RECT  3.830 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.080 0.400 ;
        RECT  1.080 -0.400 1.480 0.560 ;
        RECT  1.480 -0.400 3.530 0.400 ;
        RECT  3.530 -0.400 3.930 0.560 ;
        RECT  3.930 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.110 3.870 4.510 4.310 ;
        RECT  2.990 3.870 4.110 4.110 ;
        RECT  3.900 1.870 4.060 2.270 ;
        RECT  3.660 0.860 3.900 2.270 ;
        RECT  2.430 0.860 3.660 1.100 ;
        RECT  2.650 3.300 2.990 4.110 ;
        RECT  2.650 1.510 2.840 1.910 ;
        RECT  2.410 1.510 2.650 4.110 ;
        RECT  2.090 0.670 2.430 1.100 ;
        RECT  0.600 3.870 2.410 4.110 ;
        RECT  2.030 0.670 2.090 3.540 ;
        RECT  1.850 0.860 2.030 3.540 ;
        RECT  1.670 3.300 1.850 3.540 ;
        RECT  1.320 2.610 1.560 3.010 ;
        RECT  1.300 1.150 1.540 1.550 ;
        RECT  0.600 2.690 1.320 2.930 ;
        RECT  0.600 1.230 1.300 1.470 ;
        RECT  0.430 0.780 0.600 1.470 ;
        RECT  0.430 2.690 0.600 3.470 ;
        RECT  0.200 3.870 0.600 4.350 ;
        RECT  0.190 0.780 0.430 3.470 ;
    END
END TBUFX1

MACRO TBUFX16
    CLASS CORE ;
    FOREIGN TBUFX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFXL ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  7.330 2.910 8.790 3.890 ;
        RECT  7.160 1.140 8.790 1.940 ;
        RECT  8.790 1.140 10.350 3.890 ;
        RECT  10.350 1.140 11.630 1.940 ;
        RECT  10.350 2.910 12.380 3.890 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.700 2.250 0.950 2.650 ;
        RECT  0.950 2.240 1.210 2.660 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.330 2.070 4.820 2.470 ;
        RECT  4.820 1.830 5.080 2.470 ;
        RECT  5.080 2.070 5.310 2.470 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.760 0.170 5.440 ;
        RECT  0.170 3.560 0.570 5.440 ;
        RECT  0.570 3.760 0.580 5.440 ;
        RECT  0.580 4.630 0.680 5.440 ;
        RECT  0.680 4.640 3.820 5.440 ;
        RECT  3.820 4.280 3.830 5.440 ;
        RECT  3.830 4.080 4.230 5.440 ;
        RECT  4.230 4.280 4.240 5.440 ;
        RECT  4.240 4.640 5.300 5.440 ;
        RECT  5.300 4.210 5.310 5.440 ;
        RECT  5.310 4.010 5.710 5.440 ;
        RECT  5.710 4.210 5.720 5.440 ;
        RECT  5.720 4.640 6.710 5.440 ;
        RECT  6.710 4.370 6.720 5.440 ;
        RECT  6.720 4.170 7.120 5.440 ;
        RECT  7.120 4.370 7.130 5.440 ;
        RECT  7.130 4.640 8.110 5.440 ;
        RECT  8.110 4.370 8.120 5.440 ;
        RECT  8.120 4.170 8.520 5.440 ;
        RECT  8.520 4.370 8.530 5.440 ;
        RECT  8.530 4.640 9.680 5.440 ;
        RECT  9.680 4.370 9.690 5.440 ;
        RECT  9.690 4.170 10.090 5.440 ;
        RECT  10.090 4.370 10.100 5.440 ;
        RECT  10.100 4.640 11.220 5.440 ;
        RECT  11.220 4.370 11.230 5.440 ;
        RECT  11.230 4.170 11.630 5.440 ;
        RECT  11.630 4.370 11.640 5.440 ;
        RECT  11.640 4.640 12.620 5.440 ;
        RECT  12.620 4.370 12.630 5.440 ;
        RECT  12.630 4.170 13.030 5.440 ;
        RECT  13.030 4.370 13.040 5.440 ;
        RECT  13.040 4.640 13.200 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.330 0.400 ;
        RECT  1.330 -0.400 1.340 1.150 ;
        RECT  1.340 -0.400 1.740 1.350 ;
        RECT  1.740 -0.400 1.750 1.150 ;
        RECT  1.750 -0.400 4.240 0.400 ;
        RECT  4.240 -0.400 4.250 0.670 ;
        RECT  4.250 -0.400 4.650 0.870 ;
        RECT  4.650 -0.400 4.660 0.670 ;
        RECT  4.660 -0.400 5.580 0.400 ;
        RECT  5.580 -0.400 5.590 0.670 ;
        RECT  5.590 -0.400 5.990 0.870 ;
        RECT  5.990 -0.400 6.000 0.670 ;
        RECT  6.000 -0.400 6.560 0.400 ;
        RECT  6.560 -0.400 6.570 0.670 ;
        RECT  6.570 -0.400 6.970 0.870 ;
        RECT  6.970 -0.400 6.980 0.670 ;
        RECT  6.980 -0.400 7.820 0.400 ;
        RECT  7.820 -0.400 7.830 0.670 ;
        RECT  7.830 -0.400 8.230 0.870 ;
        RECT  8.230 -0.400 8.240 0.670 ;
        RECT  8.240 -0.400 9.160 0.400 ;
        RECT  9.160 -0.400 9.170 0.670 ;
        RECT  9.170 -0.400 9.570 0.870 ;
        RECT  9.570 -0.400 9.580 0.670 ;
        RECT  9.580 -0.400 10.500 0.400 ;
        RECT  10.500 -0.400 10.510 0.670 ;
        RECT  10.510 -0.400 10.910 0.870 ;
        RECT  10.910 -0.400 10.920 0.670 ;
        RECT  10.920 -0.400 11.840 0.400 ;
        RECT  11.840 -0.400 11.850 0.670 ;
        RECT  11.850 -0.400 12.250 0.870 ;
        RECT  12.250 -0.400 12.260 0.670 ;
        RECT  12.260 -0.400 13.200 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  7.570 2.240 8.060 2.640 ;
        RECT  6.390 2.230 7.570 2.650 ;
        RECT  6.470 1.140 6.480 1.700 ;
        RECT  6.070 1.140 6.470 1.900 ;
        RECT  6.380 2.230 6.390 2.950 ;
        RECT  6.180 2.230 6.380 3.150 ;
        RECT  5.970 2.230 6.180 3.160 ;
        RECT  6.060 1.140 6.070 1.700 ;
        RECT  4.040 1.140 6.060 1.560 ;
        RECT  3.390 2.740 5.970 3.160 ;
        RECT  4.030 1.140 4.040 1.630 ;
        RECT  3.980 1.140 4.030 1.640 ;
        RECT  3.600 0.660 3.980 1.640 ;
        RECT  2.580 0.660 3.600 1.040 ;
        RECT  3.380 2.740 3.390 3.700 ;
        RECT  3.290 2.740 3.380 4.190 ;
        RECT  3.280 1.430 3.290 4.190 ;
        RECT  2.980 1.310 3.280 4.190 ;
        RECT  2.970 1.310 2.980 3.700 ;
        RECT  1.840 3.940 2.980 4.180 ;
        RECT  2.880 1.310 2.970 3.160 ;
        RECT  2.870 1.430 2.880 3.160 ;
        RECT  2.570 0.660 2.580 1.440 ;
        RECT  2.330 0.660 2.570 3.660 ;
        RECT  2.200 0.660 2.330 1.450 ;
        RECT  2.110 1.050 2.200 1.450 ;
        RECT  1.810 1.730 2.050 3.300 ;
        RECT  1.440 3.860 1.840 4.260 ;
        RECT  0.970 1.730 1.810 1.970 ;
        RECT  1.340 3.060 1.810 3.300 ;
        RECT  0.940 3.060 1.340 3.460 ;
        RECT  0.730 1.040 0.970 1.970 ;
        RECT  0.570 1.040 0.730 1.440 ;
    END
END TBUFX16

MACRO TBUFX12
    CLASS CORE ;
    FOREIGN TBUFX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ TBUFXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER met1 ;
        RECT  6.520 3.010 8.790 3.690 ;
        RECT  6.720 1.070 8.790 1.580 ;
        RECT  8.790 1.070 10.310 3.840 ;
        RECT  10.310 1.400 10.350 3.840 ;
        END
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.340 2.280 1.880 2.750 ;
        END
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.390 2.300 5.390 2.700 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.460 5.440 ;
        RECT  1.460 4.480 1.860 5.440 ;
        RECT  1.860 4.640 4.470 5.440 ;
        RECT  4.470 3.930 4.870 5.440 ;
        RECT  4.870 4.640 6.050 5.440 ;
        RECT  6.050 3.960 6.450 5.440 ;
        RECT  6.450 4.640 7.550 5.440 ;
        RECT  7.550 4.160 7.950 5.440 ;
        RECT  7.950 4.640 9.110 5.440 ;
        RECT  9.110 4.250 9.510 5.440 ;
        RECT  9.510 4.640 10.630 5.440 ;
        RECT  10.630 4.250 11.030 5.440 ;
        RECT  11.030 4.640 11.220 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.600 0.400 ;
        RECT  1.600 -0.400 2.000 1.340 ;
        RECT  2.000 -0.400 4.460 0.400 ;
        RECT  4.460 -0.400 4.860 0.560 ;
        RECT  4.860 -0.400 5.930 0.400 ;
        RECT  5.930 -0.400 6.330 0.840 ;
        RECT  6.330 -0.400 7.370 0.400 ;
        RECT  7.370 -0.400 7.770 0.800 ;
        RECT  7.770 -0.400 8.710 0.400 ;
        RECT  8.710 -0.400 9.110 0.800 ;
        RECT  9.110 -0.400 10.050 0.400 ;
        RECT  10.050 -0.400 10.450 0.800 ;
        RECT  10.450 -0.400 11.220 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  8.290 2.320 8.430 2.560 ;
        RECT  7.530 2.320 8.290 2.680 ;
        RECT  5.960 2.440 7.530 2.680 ;
        RECT  6.060 1.890 7.240 2.130 ;
        RECT  5.820 1.320 6.060 2.130 ;
        RECT  5.720 2.440 5.960 3.210 ;
        RECT  4.280 1.320 5.820 1.560 ;
        RECT  5.590 2.970 5.720 3.210 ;
        RECT  5.190 2.970 5.590 4.250 ;
        RECT  4.150 3.300 5.190 3.540 ;
        RECT  4.120 1.230 4.280 1.560 ;
        RECT  3.820 3.180 4.150 3.580 ;
        RECT  3.960 0.670 4.120 1.560 ;
        RECT  3.880 0.670 3.960 1.470 ;
        RECT  2.770 0.670 3.880 0.910 ;
        RECT  3.580 1.850 3.820 3.580 ;
        RECT  2.460 4.110 3.800 4.350 ;
        RECT  3.320 1.850 3.580 2.090 ;
        RECT  2.650 3.340 3.580 3.580 ;
        RECT  3.320 1.230 3.520 1.470 ;
        RECT  3.080 1.230 3.320 2.090 ;
        RECT  3.060 2.600 3.300 3.000 ;
        RECT  2.770 2.600 3.060 2.840 ;
        RECT  2.530 0.670 2.770 2.840 ;
        RECT  2.250 3.340 2.650 3.760 ;
        RECT  2.360 0.890 2.530 1.290 ;
        RECT  2.220 4.000 2.460 4.350 ;
        RECT  1.090 4.000 2.220 4.240 ;
        RECT  1.230 1.680 2.170 1.920 ;
        RECT  1.070 1.020 1.230 1.920 ;
        RECT  1.070 3.420 1.090 4.240 ;
        RECT  0.850 1.020 1.070 4.240 ;
        RECT  0.830 1.020 0.850 3.820 ;
        RECT  0.690 3.420 0.830 3.820 ;
    END
END TBUFX12

MACRO SEDFFTRXL
    CLASS CORE ;
    FOREIGN SEDFFTRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.740 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.720 0.670 3.190 1.070 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.490 2.050 1.870 2.660 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.780 1.420 0.860 1.820 ;
        RECT  0.860 1.420 1.120 2.090 ;
        RECT  1.120 1.420 1.180 1.820 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  23.790 3.510 24.190 3.980 ;
        RECT  24.190 3.510 24.220 3.770 ;
        RECT  23.890 0.740 24.290 1.100 ;
        RECT  24.220 3.510 24.630 3.750 ;
        RECT  24.290 0.860 24.630 1.100 ;
        RECT  24.630 0.860 24.870 3.750 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  25.170 3.310 25.190 3.710 ;
        RECT  25.150 1.270 25.190 1.800 ;
        RECT  25.190 3.220 25.290 3.710 ;
        RECT  25.190 1.270 25.290 1.820 ;
        RECT  25.290 1.270 25.530 3.710 ;
        RECT  25.530 1.270 25.540 1.960 ;
        RECT  25.540 1.400 25.550 1.960 ;
        RECT  25.530 3.070 25.570 3.710 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.690 1.820 9.130 2.230 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.140 1.830 6.150 2.090 ;
        RECT  6.150 1.830 6.680 2.230 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  12.650 1.830 13.110 2.270 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.480 5.440 ;
        RECT  1.480 4.480 1.880 5.440 ;
        RECT  1.880 4.640 6.080 5.440 ;
        RECT  6.080 4.120 6.480 5.440 ;
        RECT  6.480 4.640 9.100 5.440 ;
        RECT  9.100 4.240 9.110 5.440 ;
        RECT  9.110 4.120 9.510 5.440 ;
        RECT  9.510 4.240 9.520 5.440 ;
        RECT  9.520 4.640 13.000 5.440 ;
        RECT  13.000 4.240 13.010 5.440 ;
        RECT  13.010 4.120 13.410 5.440 ;
        RECT  13.410 4.240 13.420 5.440 ;
        RECT  13.420 4.640 16.410 5.440 ;
        RECT  16.410 4.480 17.390 5.440 ;
        RECT  17.390 4.640 19.490 5.440 ;
        RECT  19.490 4.480 19.890 5.440 ;
        RECT  19.890 4.640 23.020 5.440 ;
        RECT  23.020 3.840 23.030 5.440 ;
        RECT  23.030 3.640 23.430 5.440 ;
        RECT  23.430 3.840 23.440 5.440 ;
        RECT  23.440 4.640 24.520 5.440 ;
        RECT  24.520 4.480 24.920 5.440 ;
        RECT  24.920 4.640 25.740 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.250 0.400 ;
        RECT  0.250 -0.400 0.650 0.560 ;
        RECT  0.650 -0.400 2.010 0.400 ;
        RECT  2.010 -0.400 2.410 0.930 ;
        RECT  2.410 -0.400 5.930 0.400 ;
        RECT  5.930 -0.400 6.330 0.560 ;
        RECT  6.330 -0.400 9.180 0.400 ;
        RECT  9.180 -0.400 9.580 1.120 ;
        RECT  9.580 -0.400 13.220 0.400 ;
        RECT  13.220 -0.400 13.620 0.560 ;
        RECT  13.620 -0.400 14.570 0.400 ;
        RECT  14.570 -0.400 14.580 1.320 ;
        RECT  14.580 -0.400 14.980 1.520 ;
        RECT  14.980 -0.400 14.990 1.320 ;
        RECT  14.990 -0.400 17.310 0.400 ;
        RECT  17.310 -0.400 17.320 1.020 ;
        RECT  17.320 -0.400 17.720 1.140 ;
        RECT  17.720 -0.400 17.730 1.020 ;
        RECT  17.730 -0.400 19.920 0.400 ;
        RECT  19.920 -0.400 20.320 1.080 ;
        RECT  20.320 -0.400 23.010 0.400 ;
        RECT  23.010 -0.400 23.410 0.560 ;
        RECT  23.410 -0.400 24.970 0.400 ;
        RECT  24.970 -0.400 25.370 0.560 ;
        RECT  25.370 -0.400 25.740 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  24.110 1.400 24.350 3.170 ;
        RECT  23.890 1.400 24.110 1.800 ;
        RECT  23.860 2.740 24.110 3.170 ;
        RECT  22.440 2.930 23.860 3.170 ;
        RECT  22.990 1.990 23.610 2.390 ;
        RECT  22.750 1.190 22.990 2.650 ;
        RECT  21.590 1.190 22.750 1.430 ;
        RECT  21.730 2.410 22.750 2.650 ;
        RECT  22.050 1.730 22.450 2.130 ;
        RECT  22.200 2.930 22.440 4.180 ;
        RECT  15.230 3.940 22.200 4.180 ;
        RECT  21.210 1.890 22.050 2.130 ;
        RECT  21.490 2.410 21.730 3.460 ;
        RECT  20.820 1.110 21.220 1.600 ;
        RECT  20.970 1.890 21.210 3.660 ;
        RECT  15.760 3.420 20.970 3.660 ;
        RECT  20.690 1.360 20.820 1.600 ;
        RECT  20.450 1.360 20.690 3.130 ;
        RECT  19.930 2.000 20.170 3.130 ;
        RECT  18.200 2.890 19.930 3.130 ;
        RECT  19.120 0.940 19.440 1.340 ;
        RECT  18.880 0.940 19.120 2.620 ;
        RECT  18.680 1.560 18.880 1.960 ;
        RECT  18.580 2.380 18.880 2.620 ;
        RECT  18.300 0.880 18.600 1.280 ;
        RECT  18.200 0.880 18.300 2.550 ;
        RECT  18.060 0.880 18.200 3.130 ;
        RECT  17.800 2.310 18.060 3.130 ;
        RECT  17.150 2.310 17.800 2.550 ;
        RECT  16.380 1.420 17.780 1.820 ;
        RECT  16.750 2.150 17.150 2.550 ;
        RECT  16.140 0.820 16.380 2.800 ;
        RECT  15.980 0.820 16.140 1.060 ;
        RECT  15.260 2.560 16.140 2.800 ;
        RECT  15.520 3.090 15.760 3.660 ;
        RECT  15.530 1.260 15.690 1.660 ;
        RECT  15.290 1.260 15.530 2.040 ;
        RECT  14.980 3.090 15.520 3.330 ;
        RECT  14.980 1.800 15.290 2.040 ;
        RECT  14.990 3.610 15.230 4.180 ;
        RECT  14.450 3.610 14.990 3.850 ;
        RECT  14.740 1.800 14.980 3.330 ;
        RECT  13.660 2.560 14.740 2.800 ;
        RECT  13.930 4.130 14.650 4.370 ;
        RECT  14.210 3.080 14.450 3.850 ;
        RECT  11.910 3.080 14.210 3.320 ;
        RECT  13.690 3.600 13.930 4.370 ;
        RECT  4.030 3.600 13.690 3.840 ;
        RECT  13.420 1.210 13.660 2.800 ;
        RECT  12.800 1.210 13.420 1.450 ;
        RECT  12.250 2.560 13.420 2.800 ;
        RECT  12.400 1.050 12.800 1.450 ;
        RECT  11.850 1.110 11.960 1.510 ;
        RECT  11.850 2.680 11.910 3.320 ;
        RECT  11.610 1.110 11.850 3.320 ;
        RECT  11.560 1.110 11.610 1.510 ;
        RECT  11.510 2.680 11.610 3.320 ;
        RECT  11.160 1.130 11.200 1.530 ;
        RECT  11.150 1.130 11.160 3.000 ;
        RECT  10.920 1.130 11.150 3.320 ;
        RECT  10.800 1.130 10.920 1.530 ;
        RECT  10.750 2.680 10.920 3.320 ;
        RECT  7.830 3.080 10.750 3.320 ;
        RECT  10.410 1.910 10.520 2.310 ;
        RECT  10.380 1.130 10.460 1.530 ;
        RECT  10.380 1.910 10.410 2.800 ;
        RECT  10.140 1.120 10.380 2.800 ;
        RECT  10.060 1.130 10.140 1.530 ;
        RECT  9.980 2.560 10.140 2.800 ;
        RECT  9.640 1.880 9.760 2.280 ;
        RECT  9.400 1.880 9.640 2.790 ;
        RECT  8.420 2.550 9.400 2.790 ;
        RECT  8.420 1.120 8.700 1.520 ;
        RECT  8.180 1.120 8.420 2.790 ;
        RECT  8.010 1.910 8.180 2.310 ;
        RECT  7.720 1.040 7.880 1.450 ;
        RECT  7.720 2.660 7.830 3.320 ;
        RECT  7.480 1.040 7.720 3.320 ;
        RECT  4.870 3.080 7.480 3.320 ;
        RECT  6.960 1.130 7.200 2.790 ;
        RECT  6.800 1.130 6.960 1.370 ;
        RECT  6.750 2.550 6.960 2.790 ;
        RECT  2.400 4.120 5.810 4.360 ;
        RECT  5.610 1.120 5.660 2.310 ;
        RECT  5.260 1.120 5.610 2.790 ;
        RECT  5.210 1.910 5.260 2.790 ;
        RECT  4.940 1.910 5.210 2.310 ;
        RECT  4.650 1.120 4.920 1.520 ;
        RECT  4.650 2.880 4.870 3.320 ;
        RECT  4.410 1.120 4.650 3.320 ;
        RECT  4.020 1.330 4.030 3.840 ;
        RECT  3.790 1.250 4.020 3.840 ;
        RECT  3.780 1.250 3.790 1.650 ;
        RECT  3.180 1.350 3.340 1.750 ;
        RECT  2.940 1.350 3.180 3.070 ;
        RECT  2.720 2.830 2.940 3.070 ;
        RECT  2.700 3.420 2.940 3.840 ;
        RECT  2.400 3.420 2.700 3.660 ;
        RECT  2.160 1.540 2.400 3.660 ;
        RECT  2.160 3.940 2.400 4.360 ;
        RECT  1.720 1.540 2.160 1.780 ;
        RECT  0.920 2.930 2.160 3.170 ;
        RECT  0.600 3.940 2.160 4.180 ;
        RECT  1.480 1.380 1.720 1.780 ;
        RECT  1.130 0.670 1.530 1.100 ;
        RECT  0.400 0.860 1.130 1.100 ;
        RECT  0.680 2.740 0.920 3.170 ;
        RECT  0.400 3.640 0.600 4.180 ;
        RECT  0.160 0.860 0.400 4.180 ;
    END
END SEDFFTRXL

MACRO SEDFFTRX4
    CLASS CORE ;
    FOREIGN SEDFFTRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SEDFFTRXL ;
    SIZE 28.380 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.720 0.710 3.190 1.110 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 2.130 1.520 2.530 ;
        RECT  1.520 2.130 1.780 2.650 ;
        RECT  1.780 2.130 1.880 2.530 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.780 1.420 0.860 1.820 ;
        RECT  0.860 1.420 1.120 2.090 ;
        RECT  1.120 1.420 1.180 1.820 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  25.620 2.750 25.850 3.150 ;
        RECT  25.840 1.150 25.850 1.660 ;
        RECT  25.850 1.150 26.240 3.150 ;
        RECT  26.240 1.260 26.250 3.150 ;
        RECT  26.250 1.260 26.290 2.660 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  27.180 1.150 27.580 1.550 ;
        RECT  27.170 2.750 27.610 4.340 ;
        RECT  27.610 2.750 27.670 3.220 ;
        RECT  27.580 1.310 27.670 1.550 ;
        RECT  27.670 1.310 27.690 3.220 ;
        RECT  27.690 1.310 27.910 3.100 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.690 1.820 9.130 2.230 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.140 1.830 6.150 2.090 ;
        RECT  6.150 1.830 6.630 2.230 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  12.710 1.880 12.740 2.280 ;
        RECT  12.740 1.830 13.110 2.280 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.840 5.440 ;
        RECT  1.840 4.480 2.240 5.440 ;
        RECT  2.240 4.640 6.080 5.440 ;
        RECT  6.080 4.120 6.480 5.440 ;
        RECT  6.480 4.640 9.040 5.440 ;
        RECT  9.040 4.240 9.050 5.440 ;
        RECT  9.050 4.120 9.450 5.440 ;
        RECT  9.450 4.240 9.460 5.440 ;
        RECT  9.460 4.640 13.000 5.440 ;
        RECT  13.000 4.240 13.010 5.440 ;
        RECT  13.010 4.120 13.410 5.440 ;
        RECT  13.410 4.240 13.420 5.440 ;
        RECT  13.420 4.640 16.410 5.440 ;
        RECT  16.410 4.480 17.390 5.440 ;
        RECT  17.390 4.640 19.550 5.440 ;
        RECT  19.550 4.480 19.950 5.440 ;
        RECT  19.950 4.640 22.990 5.440 ;
        RECT  22.740 3.680 22.990 4.080 ;
        RECT  22.990 3.680 23.390 5.440 ;
        RECT  23.390 3.680 23.640 4.080 ;
        RECT  23.390 4.640 24.850 5.440 ;
        RECT  24.850 4.120 25.250 5.440 ;
        RECT  25.250 4.640 26.310 5.440 ;
        RECT  26.310 4.040 26.710 5.440 ;
        RECT  26.710 4.640 27.890 5.440 ;
        RECT  27.890 4.010 28.130 5.440 ;
        RECT  28.130 4.640 28.380 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.250 0.400 ;
        RECT  0.250 -0.400 0.650 0.560 ;
        RECT  0.650 -0.400 2.010 0.400 ;
        RECT  2.010 -0.400 2.410 0.930 ;
        RECT  2.410 -0.400 5.830 0.400 ;
        RECT  5.830 -0.400 6.230 0.560 ;
        RECT  6.230 -0.400 9.020 0.400 ;
        RECT  9.020 -0.400 9.420 1.120 ;
        RECT  9.420 -0.400 13.060 0.400 ;
        RECT  13.060 -0.400 13.460 0.560 ;
        RECT  13.460 -0.400 14.410 0.400 ;
        RECT  14.410 -0.400 14.420 1.320 ;
        RECT  14.420 -0.400 14.820 1.520 ;
        RECT  14.820 -0.400 14.830 1.320 ;
        RECT  14.830 -0.400 17.160 0.400 ;
        RECT  17.160 -0.400 17.560 1.140 ;
        RECT  17.560 -0.400 20.490 0.400 ;
        RECT  20.490 -0.400 21.470 0.930 ;
        RECT  21.470 -0.400 23.550 0.400 ;
        RECT  23.550 -0.400 23.950 0.560 ;
        RECT  23.950 -0.400 25.200 0.400 ;
        RECT  25.200 -0.400 25.600 0.870 ;
        RECT  25.600 -0.400 26.510 0.400 ;
        RECT  26.510 -0.400 26.910 0.870 ;
        RECT  26.910 -0.400 27.800 0.400 ;
        RECT  27.800 -0.400 28.200 0.860 ;
        RECT  28.200 -0.400 28.380 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  26.930 2.220 27.430 2.460 ;
        RECT  26.690 2.220 26.930 3.730 ;
        RECT  24.360 3.490 26.690 3.730 ;
        RECT  24.520 0.710 24.760 3.170 ;
        RECT  24.360 0.710 24.520 1.110 ;
        RECT  24.360 2.930 24.520 3.170 ;
        RECT  23.960 2.930 24.360 4.320 ;
        RECT  23.850 2.290 24.250 2.690 ;
        RECT  22.380 2.930 23.960 3.170 ;
        RECT  23.630 2.290 23.850 2.650 ;
        RECT  23.390 1.190 23.630 2.650 ;
        RECT  22.380 1.190 23.390 1.430 ;
        RECT  21.730 2.410 23.390 2.650 ;
        RECT  22.710 1.730 23.110 2.130 ;
        RECT  21.210 1.890 22.710 2.130 ;
        RECT  22.140 2.930 22.380 4.180 ;
        RECT  15.170 3.940 22.140 4.180 ;
        RECT  21.490 2.410 21.730 3.460 ;
        RECT  20.690 1.370 21.350 1.610 ;
        RECT  20.970 1.890 21.210 3.660 ;
        RECT  15.700 3.420 20.970 3.660 ;
        RECT  20.450 1.370 20.690 3.140 ;
        RECT  20.370 1.370 20.450 1.610 ;
        RECT  19.930 2.000 20.170 3.140 ;
        RECT  18.280 2.900 19.930 3.140 ;
        RECT  18.960 0.950 19.280 1.350 ;
        RECT  18.720 0.950 18.960 2.620 ;
        RECT  18.580 1.560 18.720 1.960 ;
        RECT  18.560 2.380 18.720 2.620 ;
        RECT  18.280 0.860 18.440 1.260 ;
        RECT  18.040 0.860 18.280 3.140 ;
        RECT  17.800 2.310 18.040 3.140 ;
        RECT  17.240 2.310 17.800 2.550 ;
        RECT  17.360 1.420 17.760 1.820 ;
        RECT  16.410 1.500 17.360 1.740 ;
        RECT  16.840 2.150 17.240 2.550 ;
        RECT  16.170 1.500 16.410 2.800 ;
        RECT  16.160 0.810 16.220 1.050 ;
        RECT  16.160 1.500 16.170 1.740 ;
        RECT  15.260 2.560 16.170 2.800 ;
        RECT  15.920 0.810 16.160 1.740 ;
        RECT  15.820 0.810 15.920 1.050 ;
        RECT  15.460 3.090 15.700 3.660 ;
        RECT  15.370 1.350 15.530 1.750 ;
        RECT  14.980 3.090 15.460 3.330 ;
        RECT  15.130 1.350 15.370 2.040 ;
        RECT  14.930 3.610 15.170 4.180 ;
        RECT  14.980 1.800 15.130 2.040 ;
        RECT  14.740 1.800 14.980 3.330 ;
        RECT  14.450 3.610 14.930 3.850 ;
        RECT  12.380 2.560 14.740 2.800 ;
        RECT  13.930 4.130 14.650 4.370 ;
        RECT  14.210 3.080 14.450 3.850 ;
        RECT  11.850 3.080 14.210 3.320 ;
        RECT  13.690 3.600 13.930 4.370 ;
        RECT  3.920 3.600 13.690 3.840 ;
        RECT  12.380 1.050 12.640 1.450 ;
        RECT  12.140 1.050 12.380 2.800 ;
        RECT  11.690 2.680 11.850 3.320 ;
        RECT  11.690 1.110 11.800 1.510 ;
        RECT  11.450 1.110 11.690 3.320 ;
        RECT  11.400 1.110 11.450 1.510 ;
        RECT  11.000 2.680 11.090 3.320 ;
        RECT  11.000 1.120 11.040 1.520 ;
        RECT  10.760 1.120 11.000 3.320 ;
        RECT  10.640 1.120 10.760 1.520 ;
        RECT  10.690 2.680 10.760 3.320 ;
        RECT  7.850 3.080 10.690 3.320 ;
        RECT  10.410 1.910 10.480 2.310 ;
        RECT  10.320 1.910 10.410 2.800 ;
        RECT  10.080 1.120 10.320 2.800 ;
        RECT  9.900 1.120 10.080 1.520 ;
        RECT  9.920 2.560 10.080 2.800 ;
        RECT  9.640 1.880 9.760 2.280 ;
        RECT  9.400 1.880 9.640 2.790 ;
        RECT  8.370 2.550 9.400 2.790 ;
        RECT  8.460 1.130 8.540 1.530 ;
        RECT  8.370 1.120 8.460 1.530 ;
        RECT  8.130 1.120 8.370 2.790 ;
        RECT  7.950 1.910 8.130 2.310 ;
        RECT  7.670 2.660 7.850 3.320 ;
        RECT  7.670 1.040 7.720 1.450 ;
        RECT  7.430 1.040 7.670 3.320 ;
        RECT  4.760 3.080 7.430 3.320 ;
        RECT  6.910 1.130 7.150 2.800 ;
        RECT  6.640 1.130 6.910 1.370 ;
        RECT  6.690 2.560 6.910 2.800 ;
        RECT  2.790 4.120 5.810 4.360 ;
        RECT  5.560 2.040 5.610 2.790 ;
        RECT  5.210 1.050 5.560 2.790 ;
        RECT  5.160 1.050 5.210 2.440 ;
        RECT  4.720 2.040 5.160 2.440 ;
        RECT  4.440 1.050 4.820 1.490 ;
        RECT  4.440 2.880 4.760 3.320 ;
        RECT  4.420 1.050 4.440 3.320 ;
        RECT  4.200 1.250 4.420 3.320 ;
        RECT  3.920 0.730 4.000 0.970 ;
        RECT  3.680 0.730 3.920 3.840 ;
        RECT  3.600 0.730 3.680 0.970 ;
        RECT  2.400 3.400 3.400 3.640 ;
        RECT  3.180 1.390 3.340 1.790 ;
        RECT  2.940 1.390 3.180 3.060 ;
        RECT  2.720 2.820 2.940 3.060 ;
        RECT  2.550 3.940 2.790 4.360 ;
        RECT  0.840 3.940 2.550 4.180 ;
        RECT  2.160 1.540 2.400 3.640 ;
        RECT  1.720 1.540 2.160 1.780 ;
        RECT  1.160 2.930 2.160 3.170 ;
        RECT  1.480 1.380 1.720 1.780 ;
        RECT  1.130 0.670 1.530 1.100 ;
        RECT  0.920 2.740 1.160 3.170 ;
        RECT  0.500 0.860 1.130 1.100 ;
        RECT  0.500 3.640 0.840 4.180 ;
        RECT  0.260 0.860 0.500 4.180 ;
    END
END SEDFFTRX4

MACRO SEDFFTRX2
    CLASS CORE ;
    FOREIGN SEDFFTRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SEDFFTRXL ;
    SIZE 27.060 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.720 0.710 3.280 1.110 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 2.140 1.520 2.540 ;
        RECT  1.520 2.140 1.780 2.650 ;
        RECT  1.780 2.140 1.880 2.540 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.780 1.420 0.860 1.820 ;
        RECT  0.860 1.420 1.120 2.090 ;
        RECT  1.120 1.420 1.180 1.820 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  25.150 2.750 25.170 3.150 ;
        RECT  25.170 1.150 25.410 3.150 ;
        RECT  25.410 2.390 25.540 2.650 ;
        RECT  25.410 1.150 25.550 1.550 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  25.940 1.260 26.470 1.540 ;
        RECT  26.450 2.890 26.660 3.250 ;
        RECT  26.470 1.150 26.660 1.550 ;
        RECT  26.660 1.150 26.900 3.250 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.610 1.830 9.150 2.230 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.140 1.830 6.630 2.230 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  12.620 1.880 12.740 2.280 ;
        RECT  12.740 1.830 13.020 2.280 ;
        RECT  13.020 1.830 13.110 2.200 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.840 5.440 ;
        RECT  1.840 4.480 2.240 5.440 ;
        RECT  2.240 4.640 6.080 5.440 ;
        RECT  6.080 4.120 6.480 5.440 ;
        RECT  6.480 4.640 9.040 5.440 ;
        RECT  9.040 4.240 9.050 5.440 ;
        RECT  9.050 4.120 9.450 5.440 ;
        RECT  9.450 4.240 9.460 5.440 ;
        RECT  9.460 4.640 13.010 5.440 ;
        RECT  13.010 4.120 13.410 5.440 ;
        RECT  13.410 4.640 16.410 5.440 ;
        RECT  16.410 4.480 17.390 5.440 ;
        RECT  17.390 4.640 19.540 5.440 ;
        RECT  19.540 4.480 19.940 5.440 ;
        RECT  19.940 4.640 23.060 5.440 ;
        RECT  22.780 3.530 23.060 3.930 ;
        RECT  23.060 3.530 23.480 5.440 ;
        RECT  23.480 3.530 23.760 3.930 ;
        RECT  23.480 4.640 25.830 5.440 ;
        RECT  25.830 4.210 25.840 5.440 ;
        RECT  25.840 4.090 26.240 5.440 ;
        RECT  26.240 4.210 26.250 5.440 ;
        RECT  26.250 4.640 27.060 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.250 0.400 ;
        RECT  0.250 -0.400 0.650 0.560 ;
        RECT  0.650 -0.400 2.010 0.400 ;
        RECT  2.010 -0.400 2.410 0.930 ;
        RECT  2.410 -0.400 5.830 0.400 ;
        RECT  5.830 -0.400 6.230 0.560 ;
        RECT  6.230 -0.400 9.020 0.400 ;
        RECT  9.020 -0.400 9.420 1.120 ;
        RECT  9.420 -0.400 13.050 0.400 ;
        RECT  13.050 -0.400 13.450 0.560 ;
        RECT  13.450 -0.400 14.430 0.400 ;
        RECT  14.430 -0.400 14.830 1.520 ;
        RECT  14.830 -0.400 17.160 0.400 ;
        RECT  17.160 -0.400 17.560 1.140 ;
        RECT  17.560 -0.400 20.490 0.400 ;
        RECT  20.490 -0.400 21.470 0.930 ;
        RECT  21.470 -0.400 23.670 0.400 ;
        RECT  23.670 -0.400 24.070 0.560 ;
        RECT  24.070 -0.400 25.840 0.400 ;
        RECT  25.840 -0.400 25.850 0.670 ;
        RECT  25.850 -0.400 26.250 0.870 ;
        RECT  26.250 -0.400 26.260 0.670 ;
        RECT  26.260 -0.400 27.060 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  26.170 2.130 26.350 2.560 ;
        RECT  25.930 2.130 26.170 3.730 ;
        RECT  24.800 3.490 25.930 3.730 ;
        RECT  24.800 0.660 24.890 1.640 ;
        RECT  24.560 0.660 24.800 3.730 ;
        RECT  24.490 0.660 24.560 1.640 ;
        RECT  24.510 2.930 24.560 3.730 ;
        RECT  24.110 2.930 24.510 4.020 ;
        RECT  23.630 1.920 24.270 2.320 ;
        RECT  22.380 2.930 24.110 3.170 ;
        RECT  23.390 1.190 23.630 2.650 ;
        RECT  22.380 1.190 23.390 1.430 ;
        RECT  21.730 2.410 23.390 2.650 ;
        RECT  22.710 1.730 23.110 2.130 ;
        RECT  21.210 1.890 22.710 2.130 ;
        RECT  22.140 2.930 22.380 4.180 ;
        RECT  15.170 3.940 22.140 4.180 ;
        RECT  21.490 2.410 21.730 3.460 ;
        RECT  20.690 1.370 21.350 1.610 ;
        RECT  20.970 1.890 21.210 3.660 ;
        RECT  15.700 3.420 20.970 3.660 ;
        RECT  20.450 1.370 20.690 3.140 ;
        RECT  20.370 1.370 20.450 1.610 ;
        RECT  19.940 2.000 20.180 3.140 ;
        RECT  18.280 2.900 19.940 3.140 ;
        RECT  18.960 0.940 19.280 1.340 ;
        RECT  18.720 0.940 18.960 2.620 ;
        RECT  18.580 1.560 18.720 1.960 ;
        RECT  18.560 2.380 18.720 2.620 ;
        RECT  18.280 0.860 18.440 1.260 ;
        RECT  18.040 0.860 18.280 3.140 ;
        RECT  17.800 2.310 18.040 3.140 ;
        RECT  17.250 2.310 17.800 2.550 ;
        RECT  17.360 1.420 17.760 1.820 ;
        RECT  16.410 1.500 17.360 1.740 ;
        RECT  16.850 2.150 17.250 2.550 ;
        RECT  16.170 1.500 16.410 2.800 ;
        RECT  16.160 0.810 16.220 1.050 ;
        RECT  16.160 1.500 16.170 1.740 ;
        RECT  15.260 2.560 16.170 2.800 ;
        RECT  15.920 0.810 16.160 1.740 ;
        RECT  15.820 0.810 15.920 1.050 ;
        RECT  15.460 3.090 15.700 3.660 ;
        RECT  15.370 1.350 15.530 1.750 ;
        RECT  14.980 3.090 15.460 3.330 ;
        RECT  15.130 1.350 15.370 2.040 ;
        RECT  14.930 3.610 15.170 4.180 ;
        RECT  14.980 1.800 15.130 2.040 ;
        RECT  14.740 1.800 14.980 3.330 ;
        RECT  14.450 3.610 14.930 3.850 ;
        RECT  12.380 2.550 14.740 2.790 ;
        RECT  13.930 4.130 14.650 4.370 ;
        RECT  14.210 3.080 14.450 3.850 ;
        RECT  11.850 3.080 14.210 3.320 ;
        RECT  13.690 3.600 13.930 4.370 ;
        RECT  3.920 3.600 13.690 3.840 ;
        RECT  12.380 1.050 12.640 1.450 ;
        RECT  12.140 1.050 12.380 2.790 ;
        RECT  11.690 2.680 11.850 3.320 ;
        RECT  11.690 1.110 11.800 1.510 ;
        RECT  11.450 1.110 11.690 3.320 ;
        RECT  11.400 1.110 11.450 1.510 ;
        RECT  11.000 2.680 11.090 3.320 ;
        RECT  11.000 1.120 11.040 1.520 ;
        RECT  10.760 1.120 11.000 3.320 ;
        RECT  10.640 1.120 10.760 1.520 ;
        RECT  10.690 2.680 10.760 3.320 ;
        RECT  7.850 3.080 10.690 3.320 ;
        RECT  10.410 1.910 10.480 2.310 ;
        RECT  10.320 1.910 10.410 2.790 ;
        RECT  10.080 1.130 10.320 2.790 ;
        RECT  9.900 1.130 10.080 1.530 ;
        RECT  9.920 2.550 10.080 2.790 ;
        RECT  9.640 1.880 9.760 2.280 ;
        RECT  9.400 1.880 9.640 2.790 ;
        RECT  8.370 2.550 9.400 2.790 ;
        RECT  8.370 1.130 8.540 1.530 ;
        RECT  8.130 1.130 8.370 2.790 ;
        RECT  7.950 1.920 8.130 2.320 ;
        RECT  7.670 2.660 7.850 3.320 ;
        RECT  7.670 1.040 7.720 1.450 ;
        RECT  7.430 1.040 7.670 3.320 ;
        RECT  4.760 3.080 7.430 3.320 ;
        RECT  6.910 1.130 7.150 2.800 ;
        RECT  6.640 1.130 6.910 1.370 ;
        RECT  6.690 2.560 6.910 2.800 ;
        RECT  2.790 4.120 5.820 4.360 ;
        RECT  5.560 2.040 5.610 2.790 ;
        RECT  5.210 1.050 5.560 2.790 ;
        RECT  5.160 1.050 5.210 2.440 ;
        RECT  4.720 2.040 5.160 2.440 ;
        RECT  4.440 1.050 4.820 1.490 ;
        RECT  4.440 2.880 4.760 3.320 ;
        RECT  4.420 1.050 4.440 3.320 ;
        RECT  4.200 1.250 4.420 3.320 ;
        RECT  3.920 0.730 4.010 0.970 ;
        RECT  3.680 0.730 3.920 3.840 ;
        RECT  3.610 0.730 3.680 0.970 ;
        RECT  2.400 3.400 3.400 3.640 ;
        RECT  3.180 1.390 3.340 1.790 ;
        RECT  2.940 1.390 3.180 3.060 ;
        RECT  2.720 2.820 2.940 3.060 ;
        RECT  2.550 3.940 2.790 4.360 ;
        RECT  0.840 3.940 2.550 4.180 ;
        RECT  2.160 1.540 2.400 3.640 ;
        RECT  1.720 1.540 2.160 1.780 ;
        RECT  1.160 2.930 2.160 3.170 ;
        RECT  1.480 1.380 1.720 1.780 ;
        RECT  1.130 0.670 1.530 1.100 ;
        RECT  0.920 2.740 1.160 3.170 ;
        RECT  0.500 0.860 1.130 1.100 ;
        RECT  0.500 3.640 0.840 4.180 ;
        RECT  0.260 0.860 0.500 4.180 ;
    END
END SEDFFTRX2

MACRO SEDFFTRX1
    CLASS CORE ;
    FOREIGN SEDFFTRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SEDFFTRXL ;
    SIZE 27.060 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.640 0.710 3.190 1.110 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 2.130 1.520 2.530 ;
        RECT  1.520 2.130 1.780 2.650 ;
        RECT  1.780 2.130 1.880 2.530 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.740 1.410 0.770 1.810 ;
        RECT  0.770 1.410 0.860 1.820 ;
        RECT  0.860 1.410 1.120 2.090 ;
        RECT  1.120 1.410 1.140 1.820 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  25.070 1.400 25.190 1.800 ;
        RECT  24.850 3.120 25.250 3.520 ;
        RECT  25.250 3.120 25.290 3.360 ;
        RECT  25.280 2.390 25.290 2.650 ;
        RECT  25.190 1.400 25.290 1.820 ;
        RECT  25.290 1.400 25.530 3.360 ;
        RECT  25.530 2.390 25.540 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  25.940 1.270 26.290 1.530 ;
        RECT  26.290 1.270 26.490 1.540 ;
        RECT  26.490 1.270 26.610 1.670 ;
        RECT  26.490 2.880 26.650 3.280 ;
        RECT  26.610 1.270 26.650 1.840 ;
        RECT  26.650 1.270 26.890 3.280 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.610 1.830 9.130 2.230 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.140 1.830 6.630 2.230 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  12.710 1.880 12.740 2.280 ;
        RECT  12.740 1.830 13.110 2.280 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.840 5.440 ;
        RECT  1.840 4.480 2.240 5.440 ;
        RECT  2.240 4.640 6.080 5.440 ;
        RECT  6.080 4.120 6.480 5.440 ;
        RECT  6.480 4.640 9.050 5.440 ;
        RECT  9.050 4.120 9.450 5.440 ;
        RECT  9.450 4.640 13.010 5.440 ;
        RECT  13.010 4.120 13.410 5.440 ;
        RECT  13.410 4.640 16.410 5.440 ;
        RECT  16.410 4.480 17.390 5.440 ;
        RECT  17.390 4.640 19.540 5.440 ;
        RECT  19.540 4.480 19.940 5.440 ;
        RECT  19.940 4.640 23.060 5.440 ;
        RECT  22.780 3.530 23.060 3.930 ;
        RECT  23.060 3.530 23.480 5.440 ;
        RECT  23.480 3.530 23.760 3.930 ;
        RECT  23.480 4.640 25.670 5.440 ;
        RECT  25.670 4.480 26.070 5.440 ;
        RECT  26.070 4.640 27.060 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.250 0.400 ;
        RECT  0.250 -0.400 0.650 0.560 ;
        RECT  0.650 -0.400 2.000 0.400 ;
        RECT  2.000 -0.400 2.400 0.930 ;
        RECT  2.400 -0.400 5.830 0.400 ;
        RECT  5.830 -0.400 6.230 0.560 ;
        RECT  6.230 -0.400 9.020 0.400 ;
        RECT  9.020 -0.400 9.420 1.120 ;
        RECT  9.420 -0.400 13.050 0.400 ;
        RECT  13.050 -0.400 13.450 0.560 ;
        RECT  13.450 -0.400 14.430 0.400 ;
        RECT  14.430 -0.400 14.830 1.520 ;
        RECT  14.830 -0.400 17.160 0.400 ;
        RECT  17.160 -0.400 17.560 1.140 ;
        RECT  17.560 -0.400 20.490 0.400 ;
        RECT  20.490 -0.400 21.470 0.930 ;
        RECT  21.470 -0.400 23.670 0.400 ;
        RECT  23.670 -0.400 24.070 0.560 ;
        RECT  24.070 -0.400 25.730 0.400 ;
        RECT  25.730 -0.400 26.130 0.560 ;
        RECT  26.130 -0.400 27.060 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  26.200 2.180 26.350 2.580 ;
        RECT  25.960 2.180 26.200 4.040 ;
        RECT  24.510 3.800 25.960 4.040 ;
        RECT  24.790 0.720 24.890 0.960 ;
        RECT  24.550 0.720 24.790 2.840 ;
        RECT  24.490 0.720 24.550 0.960 ;
        RECT  24.510 2.600 24.550 2.840 ;
        RECT  24.270 2.600 24.510 4.040 ;
        RECT  24.110 2.930 24.270 3.730 ;
        RECT  23.630 1.920 24.260 2.320 ;
        RECT  22.380 2.930 24.110 3.170 ;
        RECT  23.390 1.190 23.630 2.650 ;
        RECT  22.380 1.190 23.390 1.430 ;
        RECT  21.730 2.410 23.390 2.650 ;
        RECT  22.710 1.730 23.110 2.130 ;
        RECT  21.210 1.890 22.710 2.130 ;
        RECT  22.140 2.930 22.380 4.180 ;
        RECT  15.170 3.940 22.140 4.180 ;
        RECT  21.490 2.410 21.730 3.460 ;
        RECT  20.690 1.370 21.350 1.610 ;
        RECT  20.970 1.890 21.210 3.660 ;
        RECT  15.700 3.420 20.970 3.660 ;
        RECT  20.450 1.370 20.690 3.140 ;
        RECT  20.370 1.370 20.450 1.610 ;
        RECT  19.930 2.000 20.170 3.140 ;
        RECT  18.280 2.900 19.930 3.140 ;
        RECT  18.960 0.950 19.280 1.350 ;
        RECT  18.720 0.950 18.960 2.620 ;
        RECT  18.580 1.560 18.720 1.960 ;
        RECT  18.560 2.380 18.720 2.620 ;
        RECT  18.280 0.900 18.440 1.300 ;
        RECT  18.040 0.900 18.280 3.140 ;
        RECT  17.800 2.310 18.040 3.140 ;
        RECT  17.240 2.310 17.800 2.550 ;
        RECT  17.360 1.420 17.760 1.820 ;
        RECT  16.410 1.500 17.360 1.740 ;
        RECT  16.840 2.150 17.240 2.550 ;
        RECT  16.170 1.500 16.410 2.800 ;
        RECT  16.160 0.810 16.220 1.050 ;
        RECT  16.160 1.500 16.170 1.740 ;
        RECT  15.260 2.560 16.170 2.800 ;
        RECT  15.920 0.810 16.160 1.740 ;
        RECT  15.820 0.810 15.920 1.050 ;
        RECT  15.460 3.090 15.700 3.660 ;
        RECT  15.370 1.350 15.530 1.750 ;
        RECT  14.980 3.090 15.460 3.330 ;
        RECT  15.130 1.350 15.370 2.040 ;
        RECT  14.930 3.610 15.170 4.180 ;
        RECT  14.980 1.800 15.130 2.040 ;
        RECT  14.740 1.800 14.980 3.330 ;
        RECT  14.450 3.610 14.930 3.850 ;
        RECT  12.380 2.560 14.740 2.800 ;
        RECT  13.930 4.090 14.650 4.330 ;
        RECT  14.210 3.080 14.450 3.850 ;
        RECT  11.850 3.080 14.210 3.320 ;
        RECT  13.690 3.600 13.930 4.330 ;
        RECT  3.920 3.600 13.690 3.840 ;
        RECT  12.380 1.050 12.640 1.450 ;
        RECT  12.140 1.050 12.380 2.800 ;
        RECT  11.690 2.680 11.850 3.320 ;
        RECT  11.690 1.110 11.800 1.510 ;
        RECT  11.450 1.110 11.690 3.320 ;
        RECT  11.400 1.110 11.450 1.510 ;
        RECT  11.000 2.680 11.090 3.320 ;
        RECT  11.000 1.120 11.040 1.520 ;
        RECT  10.760 1.120 11.000 3.320 ;
        RECT  10.640 1.120 10.760 1.520 ;
        RECT  10.690 2.680 10.760 3.320 ;
        RECT  7.850 3.080 10.690 3.320 ;
        RECT  10.410 1.910 10.480 2.310 ;
        RECT  10.320 1.910 10.410 2.800 ;
        RECT  10.080 1.130 10.320 2.800 ;
        RECT  9.900 1.130 10.080 1.530 ;
        RECT  9.920 2.560 10.080 2.800 ;
        RECT  9.640 1.880 9.760 2.280 ;
        RECT  9.400 1.880 9.640 2.790 ;
        RECT  8.370 2.550 9.400 2.790 ;
        RECT  8.370 1.120 8.540 1.520 ;
        RECT  8.130 1.120 8.370 2.790 ;
        RECT  7.950 1.920 8.130 2.320 ;
        RECT  7.670 2.660 7.850 3.320 ;
        RECT  7.670 1.040 7.720 1.450 ;
        RECT  7.430 1.040 7.670 3.320 ;
        RECT  4.760 3.080 7.430 3.320 ;
        RECT  6.910 1.130 7.150 2.800 ;
        RECT  6.640 1.130 6.910 1.370 ;
        RECT  6.690 2.560 6.910 2.800 ;
        RECT  2.790 4.120 5.810 4.360 ;
        RECT  5.560 2.030 5.610 2.800 ;
        RECT  5.210 1.050 5.560 2.800 ;
        RECT  5.160 1.050 5.210 2.430 ;
        RECT  4.680 2.030 5.160 2.430 ;
        RECT  4.440 1.050 4.800 1.490 ;
        RECT  4.440 2.880 4.760 3.320 ;
        RECT  4.400 1.050 4.440 3.320 ;
        RECT  4.200 1.250 4.400 3.320 ;
        RECT  3.920 0.750 4.010 0.990 ;
        RECT  3.680 0.750 3.920 3.840 ;
        RECT  3.610 0.750 3.680 0.990 ;
        RECT  2.400 3.400 3.400 3.640 ;
        RECT  3.180 1.390 3.340 1.790 ;
        RECT  2.940 1.390 3.180 3.060 ;
        RECT  2.720 2.820 2.940 3.060 ;
        RECT  2.550 3.940 2.790 4.360 ;
        RECT  0.840 3.940 2.550 4.180 ;
        RECT  2.160 1.540 2.400 3.640 ;
        RECT  1.720 1.540 2.160 1.780 ;
        RECT  1.160 2.930 2.160 3.170 ;
        RECT  1.480 1.380 1.720 1.780 ;
        RECT  1.130 0.670 1.530 1.100 ;
        RECT  0.920 2.740 1.160 3.170 ;
        RECT  0.500 0.860 1.130 1.100 ;
        RECT  0.500 3.640 0.840 4.180 ;
        RECT  0.260 0.860 0.500 4.180 ;
    END
END SEDFFTRX1

MACRO SEDFFHQXL
    CLASS CORE ;
    FOREIGN SEDFFHQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.780 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.530 0.720 1.830 1.030 ;
        RECT  1.830 0.710 1.930 1.030 ;
        RECT  1.930 0.710 2.440 0.980 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.710 2.010 0.860 2.640 ;
        RECT  0.860 2.010 1.120 2.650 ;
        RECT  1.120 2.010 1.160 2.640 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.180 0.700 21.230 1.100 ;
        RECT  21.000 3.040 21.330 3.440 ;
        RECT  21.320 1.830 21.330 2.090 ;
        RECT  21.230 0.700 21.330 1.260 ;
        RECT  21.330 0.700 21.400 3.440 ;
        RECT  21.400 0.700 21.570 3.280 ;
        RECT  21.570 1.830 21.580 2.090 ;
        RECT  21.570 0.700 21.580 1.390 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.640 1.650 8.120 1.890 ;
        RECT  8.120 1.650 8.370 2.090 ;
        RECT  8.370 1.830 8.380 2.090 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.820 1.830 4.960 2.090 ;
        RECT  4.960 1.810 5.360 2.210 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  10.740 1.740 11.260 2.140 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.960 5.440 ;
        RECT  0.960 4.480 1.360 5.440 ;
        RECT  1.360 4.640 4.870 5.440 ;
        RECT  4.870 4.480 5.270 5.440 ;
        RECT  5.270 4.640 7.880 5.440 ;
        RECT  7.880 4.480 8.280 5.440 ;
        RECT  8.280 4.640 11.200 5.440 ;
        RECT  11.200 3.840 11.600 5.440 ;
        RECT  11.600 4.640 14.120 5.440 ;
        RECT  14.120 4.480 15.100 5.440 ;
        RECT  15.100 4.640 19.320 5.440 ;
        RECT  19.320 4.480 19.720 5.440 ;
        RECT  19.720 4.640 20.900 5.440 ;
        RECT  20.900 4.480 21.300 5.440 ;
        RECT  21.300 4.640 21.780 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 4.590 0.400 ;
        RECT  4.590 -0.400 4.990 0.560 ;
        RECT  4.990 -0.400 7.780 0.400 ;
        RECT  7.780 -0.400 8.180 0.560 ;
        RECT  8.180 -0.400 11.380 0.400 ;
        RECT  11.380 -0.400 11.780 0.560 ;
        RECT  11.780 -0.400 14.040 0.400 ;
        RECT  14.040 -0.400 14.440 0.910 ;
        RECT  14.440 -0.400 16.660 0.400 ;
        RECT  16.660 -0.400 16.900 1.140 ;
        RECT  16.900 -0.400 19.560 0.400 ;
        RECT  19.560 -0.400 19.800 1.820 ;
        RECT  19.800 -0.400 20.320 0.400 ;
        RECT  20.320 -0.400 20.720 0.560 ;
        RECT  20.720 -0.400 21.780 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  20.660 1.420 20.740 1.820 ;
        RECT  20.480 1.420 20.660 3.140 ;
        RECT  20.420 1.420 20.480 3.800 ;
        RECT  20.340 1.420 20.420 1.820 ;
        RECT  20.260 2.740 20.420 3.800 ;
        RECT  20.240 2.900 20.260 3.800 ;
        RECT  19.980 3.400 20.240 3.800 ;
        RECT  19.230 2.060 20.000 2.460 ;
        RECT  19.300 3.480 19.980 3.720 ;
        RECT  19.060 2.860 19.300 3.720 ;
        RECT  18.990 0.690 19.230 2.580 ;
        RECT  19.000 3.480 19.060 3.720 ;
        RECT  18.760 3.480 19.000 4.400 ;
        RECT  18.160 0.690 18.990 0.930 ;
        RECT  18.320 2.340 18.990 2.580 ;
        RECT  15.600 4.160 18.760 4.400 ;
        RECT  18.590 1.320 18.750 1.560 ;
        RECT  18.350 1.320 18.590 2.100 ;
        RECT  17.840 1.860 18.350 2.100 ;
        RECT  18.080 2.340 18.320 3.340 ;
        RECT  17.380 0.770 17.840 1.010 ;
        RECT  17.600 1.860 17.840 3.920 ;
        RECT  16.140 3.680 17.600 3.920 ;
        RECT  17.360 0.770 17.380 1.620 ;
        RECT  17.140 0.770 17.360 3.340 ;
        RECT  17.120 1.380 17.140 3.340 ;
        RECT  16.640 1.970 16.880 2.370 ;
        RECT  16.470 2.130 16.640 2.370 ;
        RECT  16.230 2.130 16.470 3.120 ;
        RECT  15.220 2.880 16.230 3.120 ;
        RECT  15.900 3.420 16.140 3.920 ;
        RECT  15.720 0.820 16.120 1.220 ;
        RECT  15.700 2.400 15.920 2.640 ;
        RECT  12.570 3.420 15.900 3.660 ;
        RECT  15.700 0.980 15.720 1.220 ;
        RECT  15.460 0.980 15.700 2.640 ;
        RECT  15.360 3.940 15.600 4.400 ;
        RECT  12.080 3.940 15.360 4.180 ;
        RECT  14.980 0.930 15.220 3.120 ;
        RECT  14.220 2.880 14.980 3.120 ;
        RECT  14.320 1.150 14.560 1.800 ;
        RECT  13.240 1.150 14.320 1.390 ;
        RECT  13.980 2.240 14.220 3.120 ;
        RECT  13.820 2.240 13.980 2.640 ;
        RECT  13.000 0.910 13.240 3.140 ;
        RECT  12.710 0.910 13.000 1.150 ;
        RECT  12.870 2.730 13.000 3.140 ;
        RECT  12.570 1.430 12.720 1.830 ;
        RECT  12.330 1.430 12.570 3.660 ;
        RECT  11.940 1.430 12.330 1.670 ;
        RECT  10.700 2.800 12.330 3.040 ;
        RECT  11.840 3.320 12.080 4.180 ;
        RECT  11.700 1.220 11.940 1.670 ;
        RECT  10.360 3.320 11.840 3.560 ;
        RECT  11.110 1.220 11.700 1.460 ;
        RECT  10.710 1.060 11.110 1.460 ;
        RECT  10.460 3.880 10.860 4.360 ;
        RECT  8.800 4.120 10.460 4.360 ;
        RECT  10.280 1.330 10.360 1.730 ;
        RECT  10.280 3.140 10.360 3.560 ;
        RECT  10.040 1.330 10.280 3.560 ;
        RECT  9.960 1.330 10.040 1.730 ;
        RECT  9.960 3.140 10.040 3.560 ;
        RECT  9.440 1.330 9.680 3.840 ;
        RECT  9.280 1.330 9.440 1.730 ;
        RECT  9.200 3.410 9.440 3.840 ;
        RECT  6.700 3.410 9.200 3.650 ;
        RECT  9.000 2.200 9.160 3.100 ;
        RECT  9.000 0.670 9.060 0.910 ;
        RECT  8.920 0.670 9.000 3.100 ;
        RECT  8.760 0.670 8.920 2.520 ;
        RECT  8.700 2.860 8.920 3.100 ;
        RECT  8.560 3.940 8.800 4.360 ;
        RECT  8.660 0.670 8.760 1.100 ;
        RECT  7.070 0.860 8.660 1.100 ;
        RECT  2.920 3.940 8.560 4.180 ;
        RECT  7.460 2.370 8.480 2.610 ;
        RECT  7.060 2.370 7.460 3.130 ;
        RECT  7.060 1.380 7.360 1.620 ;
        RECT  6.830 0.670 7.070 1.100 ;
        RECT  6.820 1.380 7.060 2.610 ;
        RECT  6.020 0.670 6.830 0.910 ;
        RECT  6.740 2.180 6.820 2.610 ;
        RECT  6.460 2.960 6.700 3.650 ;
        RECT  6.460 1.230 6.540 1.630 ;
        RECT  6.220 1.230 6.460 3.650 ;
        RECT  3.650 3.410 6.220 3.650 ;
        RECT  5.700 1.280 5.940 3.120 ;
        RECT  5.460 1.280 5.700 1.520 ;
        RECT  5.540 2.880 5.700 3.120 ;
        RECT  4.190 2.890 4.400 3.130 ;
        RECT  4.190 1.590 4.200 2.530 ;
        RECT  3.950 1.390 4.190 3.130 ;
        RECT  3.790 1.390 3.950 2.530 ;
        RECT  3.780 1.590 3.790 2.530 ;
        RECT  3.730 2.120 3.780 2.520 ;
        RECT  3.450 0.680 3.750 0.920 ;
        RECT  3.450 3.050 3.650 3.650 ;
        RECT  3.210 0.680 3.450 3.650 ;
        RECT  2.810 1.400 2.930 1.800 ;
        RECT  2.810 2.990 2.920 4.180 ;
        RECT  2.680 1.400 2.810 4.180 ;
        RECT  2.570 1.400 2.680 3.390 ;
        RECT  2.530 1.400 2.570 1.800 ;
        RECT  2.490 2.990 2.570 3.390 ;
        RECT  2.000 3.940 2.400 4.340 ;
        RECT  2.040 1.400 2.170 1.800 ;
        RECT  2.040 2.980 2.120 3.380 ;
        RECT  1.800 1.400 2.040 3.380 ;
        RECT  0.560 3.940 2.000 4.180 ;
        RECT  1.770 1.400 1.800 1.800 ;
        RECT  1.720 2.980 1.800 3.380 ;
        RECT  0.400 1.330 0.570 1.730 ;
        RECT  0.400 2.980 0.560 4.180 ;
        RECT  0.320 1.330 0.400 4.180 ;
        RECT  0.160 1.330 0.320 3.390 ;
    END
END SEDFFHQXL

MACRO SEDFFHQX4
    CLASS CORE ;
    FOREIGN SEDFFHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SEDFFHQXL ;
    SIZE 27.060 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.550 0.720 1.880 1.030 ;
        RECT  1.880 0.720 2.180 1.040 ;
        RECT  2.180 0.710 2.440 1.040 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.670 2.020 1.120 2.650 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  25.860 1.390 26.060 1.790 ;
        RECT  25.850 2.850 26.290 4.340 ;
        RECT  26.290 2.850 26.450 3.270 ;
        RECT  26.060 1.380 26.450 1.800 ;
        RECT  26.450 1.380 26.870 3.270 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.560 1.780 8.120 2.020 ;
        RECT  8.120 1.780 8.380 2.090 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.820 1.830 4.970 2.090 ;
        RECT  4.970 1.750 5.370 2.150 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  10.760 1.740 11.150 2.100 ;
        RECT  11.150 1.740 11.160 2.150 ;
        RECT  11.160 1.750 11.550 2.150 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.940 5.440 ;
        RECT  0.940 4.480 1.340 5.440 ;
        RECT  1.340 4.640 4.980 5.440 ;
        RECT  4.980 4.480 5.380 5.440 ;
        RECT  5.380 4.640 7.880 5.440 ;
        RECT  7.880 4.480 8.280 5.440 ;
        RECT  8.280 4.640 11.350 5.440 ;
        RECT  11.350 4.480 11.750 5.440 ;
        RECT  11.750 4.640 13.220 5.440 ;
        RECT  13.220 4.480 14.200 5.440 ;
        RECT  14.200 4.640 22.960 5.440 ;
        RECT  22.960 4.480 23.940 5.440 ;
        RECT  23.940 4.640 25.150 5.440 ;
        RECT  25.150 4.110 25.570 5.440 ;
        RECT  25.570 4.640 26.570 5.440 ;
        RECT  26.570 4.120 26.810 5.440 ;
        RECT  26.810 4.640 27.060 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.850 0.400 ;
        RECT  0.850 -0.400 1.250 0.560 ;
        RECT  1.250 -0.400 4.420 0.400 ;
        RECT  4.420 -0.400 4.820 0.560 ;
        RECT  4.820 -0.400 7.580 0.400 ;
        RECT  7.580 -0.400 7.980 0.560 ;
        RECT  7.980 -0.400 11.620 0.400 ;
        RECT  11.620 -0.400 12.020 0.560 ;
        RECT  12.020 -0.400 14.280 0.400 ;
        RECT  14.280 -0.400 14.680 1.120 ;
        RECT  14.680 -0.400 17.620 0.400 ;
        RECT  17.620 -0.400 18.020 1.520 ;
        RECT  18.020 -0.400 19.130 0.400 ;
        RECT  19.130 -0.400 19.140 1.190 ;
        RECT  19.140 -0.400 19.540 1.390 ;
        RECT  19.540 -0.400 19.550 1.190 ;
        RECT  19.550 -0.400 23.600 0.400 ;
        RECT  23.600 -0.400 24.000 0.560 ;
        RECT  24.000 -0.400 25.220 0.400 ;
        RECT  25.220 -0.400 25.620 1.100 ;
        RECT  25.620 -0.400 26.490 0.400 ;
        RECT  26.490 -0.400 26.890 1.110 ;
        RECT  26.890 -0.400 27.060 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  25.560 2.070 26.180 2.470 ;
        RECT  25.320 1.410 25.560 3.550 ;
        RECT  24.800 1.410 25.320 1.650 ;
        RECT  24.750 3.310 25.320 3.550 ;
        RECT  23.920 2.240 25.050 2.640 ;
        RECT  24.400 1.250 24.800 1.650 ;
        RECT  24.330 3.310 24.750 3.880 ;
        RECT  22.850 3.640 24.330 3.880 ;
        RECT  23.680 0.860 23.920 3.270 ;
        RECT  22.650 0.860 23.680 1.100 ;
        RECT  22.090 3.030 23.680 3.270 ;
        RECT  23.140 1.380 23.380 2.670 ;
        RECT  21.830 1.380 23.140 1.620 ;
        RECT  21.330 2.430 23.140 2.670 ;
        RECT  20.670 1.900 22.850 2.140 ;
        RECT  22.690 3.640 22.850 4.040 ;
        RECT  22.450 3.640 22.690 4.400 ;
        RECT  22.250 0.700 22.650 1.100 ;
        RECT  14.710 4.160 22.450 4.400 ;
        RECT  21.070 0.700 22.250 0.940 ;
        RECT  21.850 3.030 22.090 3.850 ;
        RECT  21.690 3.350 21.850 3.850 ;
        RECT  21.430 1.240 21.830 1.620 ;
        RECT  20.490 3.610 21.690 3.850 ;
        RECT  20.310 1.380 21.430 1.620 ;
        RECT  21.090 2.430 21.330 3.280 ;
        RECT  20.930 2.880 21.090 3.280 ;
        RECT  20.670 0.700 21.070 1.100 ;
        RECT  20.430 1.900 20.670 2.660 ;
        RECT  20.250 3.440 20.490 3.850 ;
        RECT  20.250 2.260 20.430 2.660 ;
        RECT  20.150 1.130 20.310 1.620 ;
        RECT  19.970 2.420 20.250 2.660 ;
        RECT  19.910 1.130 20.150 1.920 ;
        RECT  19.730 2.420 19.970 3.920 ;
        RECT  18.780 1.680 19.910 1.920 ;
        RECT  15.350 3.680 19.730 3.920 ;
        RECT  18.620 2.930 19.450 3.330 ;
        RECT  18.620 1.130 18.780 1.920 ;
        RECT  18.380 1.130 18.620 3.330 ;
        RECT  17.690 2.930 18.380 3.330 ;
        RECT  17.700 2.130 18.100 2.530 ;
        RECT  17.160 2.290 17.700 2.530 ;
        RECT  16.640 1.120 17.260 1.520 ;
        RECT  16.920 2.290 17.160 3.440 ;
        RECT  15.870 3.200 16.920 3.440 ;
        RECT  16.400 0.640 16.640 2.960 ;
        RECT  15.680 0.640 16.400 0.880 ;
        RECT  16.180 2.720 16.400 2.960 ;
        RECT  15.630 1.210 15.870 3.440 ;
        RECT  15.110 1.210 15.630 1.450 ;
        RECT  14.310 2.900 15.630 3.140 ;
        RECT  15.110 3.420 15.350 3.920 ;
        RECT  14.830 1.940 15.230 2.340 ;
        RECT  13.150 3.420 15.110 3.660 ;
        RECT  14.590 1.360 14.830 2.340 ;
        RECT  14.470 3.940 14.710 4.400 ;
        RECT  13.660 1.360 14.590 1.600 ;
        RECT  12.630 3.940 14.470 4.180 ;
        RECT  14.070 1.850 14.310 3.140 ;
        RECT  13.420 1.020 13.660 3.140 ;
        RECT  12.950 1.020 13.420 1.260 ;
        RECT  12.960 2.800 13.150 3.660 ;
        RECT  12.910 1.600 12.960 3.660 ;
        RECT  12.720 1.600 12.910 3.040 ;
        RECT  12.380 1.600 12.720 1.840 ;
        RECT  10.930 2.800 12.720 3.040 ;
        RECT  12.390 3.440 12.630 4.180 ;
        RECT  10.430 3.440 12.390 3.680 ;
        RECT  12.140 1.100 12.380 1.840 ;
        RECT  11.210 1.100 12.140 1.340 ;
        RECT  10.960 3.920 12.110 4.160 ;
        RECT  10.810 0.940 11.210 1.340 ;
        RECT  10.720 3.920 10.960 4.360 ;
        RECT  10.530 2.720 10.930 3.120 ;
        RECT  8.980 4.120 10.720 4.360 ;
        RECT  10.230 0.920 10.470 1.320 ;
        RECT  10.230 3.440 10.430 3.880 ;
        RECT  9.990 0.920 10.230 3.880 ;
        RECT  9.470 0.920 9.710 3.820 ;
        RECT  9.270 0.920 9.470 1.320 ;
        RECT  9.270 3.360 9.470 3.820 ;
        RECT  6.750 3.360 9.270 3.600 ;
        RECT  8.980 2.200 9.180 3.080 ;
        RECT  8.740 0.740 8.980 3.080 ;
        RECT  8.740 3.880 8.980 4.360 ;
        RECT  8.440 0.740 8.740 1.040 ;
        RECT  2.960 3.880 8.740 4.120 ;
        RECT  7.150 0.800 8.440 1.040 ;
        RECT  8.200 2.440 8.440 2.840 ;
        RECT  7.490 2.600 8.200 2.840 ;
        RECT  7.330 2.600 7.490 3.120 ;
        RECT  7.150 2.350 7.330 3.120 ;
        RECT  7.150 1.380 7.320 1.620 ;
        RECT  6.910 0.680 7.150 1.040 ;
        RECT  7.090 1.380 7.150 3.120 ;
        RECT  6.910 1.380 7.090 2.590 ;
        RECT  5.900 0.680 6.910 0.920 ;
        RECT  6.790 2.190 6.910 2.590 ;
        RECT  6.510 3.040 6.750 3.600 ;
        RECT  6.510 1.230 6.560 1.470 ;
        RECT  6.270 1.230 6.510 3.600 ;
        RECT  6.160 1.230 6.270 1.470 ;
        RECT  3.680 3.360 6.270 3.600 ;
        RECT  5.890 2.840 5.990 3.080 ;
        RECT  5.650 1.230 5.890 3.080 ;
        RECT  5.290 1.230 5.650 1.470 ;
        RECT  5.590 2.840 5.650 3.080 ;
        RECT  4.430 2.830 4.510 3.070 ;
        RECT  4.190 2.290 4.430 3.070 ;
        RECT  4.000 2.290 4.190 2.530 ;
        RECT  4.110 2.830 4.190 3.070 ;
        RECT  3.760 1.290 4.000 2.530 ;
        RECT  3.520 3.180 3.680 3.600 ;
        RECT  3.520 0.640 3.550 0.880 ;
        RECT  3.280 0.640 3.520 3.600 ;
        RECT  3.150 0.640 3.280 0.880 ;
        RECT  2.720 1.330 2.960 4.120 ;
        RECT  2.640 1.330 2.720 1.740 ;
        RECT  2.560 2.980 2.720 3.380 ;
        RECT  2.000 3.630 2.400 4.030 ;
        RECT  2.020 1.340 2.100 1.740 ;
        RECT  2.020 2.980 2.100 3.380 ;
        RECT  1.780 1.340 2.020 3.380 ;
        RECT  0.580 3.630 2.000 3.870 ;
        RECT  1.700 1.340 1.780 1.740 ;
        RECT  1.700 2.980 1.780 3.380 ;
        RECT  0.400 1.340 0.580 1.740 ;
        RECT  0.400 2.980 0.580 3.870 ;
        RECT  0.340 1.340 0.400 3.870 ;
        RECT  0.160 1.340 0.340 3.390 ;
    END
END SEDFFHQX4

MACRO SEDFFHQX2
    CLASS CORE ;
    FOREIGN SEDFFHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SEDFFHQXL ;
    SIZE 24.420 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.550 0.700 1.950 1.030 ;
        RECT  1.950 0.700 2.440 0.980 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.670 2.020 1.120 2.650 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  23.300 1.270 23.310 1.530 ;
        RECT  23.310 1.250 23.850 1.560 ;
        RECT  23.850 2.860 23.930 3.260 ;
        RECT  23.850 1.250 23.930 1.650 ;
        RECT  23.930 1.250 24.170 3.260 ;
        RECT  24.170 2.400 24.250 3.260 ;
        RECT  24.170 1.250 24.250 1.960 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.590 1.780 8.120 2.020 ;
        RECT  8.120 1.780 8.370 2.090 ;
        RECT  8.370 1.830 8.380 2.090 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.820 1.830 4.980 2.090 ;
        RECT  4.980 1.750 5.380 2.150 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  10.760 1.710 11.160 2.130 ;
        RECT  11.160 1.720 11.550 2.120 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.940 5.440 ;
        RECT  0.940 4.480 1.340 5.440 ;
        RECT  1.340 4.640 4.980 5.440 ;
        RECT  4.980 4.480 5.380 5.440 ;
        RECT  5.380 4.640 7.880 5.440 ;
        RECT  7.880 4.480 8.280 5.440 ;
        RECT  8.280 4.640 11.670 5.440 ;
        RECT  11.670 3.990 11.910 5.440 ;
        RECT  11.910 4.640 13.640 5.440 ;
        RECT  13.640 4.480 14.040 5.440 ;
        RECT  14.040 4.640 21.630 5.440 ;
        RECT  21.630 4.480 22.090 5.440 ;
        RECT  22.090 4.640 23.240 5.440 ;
        RECT  23.240 4.120 23.640 5.440 ;
        RECT  23.640 4.640 24.420 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.860 0.400 ;
        RECT  0.860 -0.400 1.260 0.560 ;
        RECT  1.260 -0.400 4.420 0.400 ;
        RECT  4.420 -0.400 4.820 0.560 ;
        RECT  4.820 -0.400 7.570 0.400 ;
        RECT  7.570 -0.400 7.970 0.560 ;
        RECT  7.970 -0.400 11.620 0.400 ;
        RECT  11.620 -0.400 12.020 0.560 ;
        RECT  12.020 -0.400 14.250 0.400 ;
        RECT  14.250 -0.400 14.650 1.090 ;
        RECT  14.650 -0.400 16.830 0.400 ;
        RECT  16.830 -0.400 17.230 1.540 ;
        RECT  17.230 -0.400 18.440 0.400 ;
        RECT  18.440 -0.400 18.680 1.650 ;
        RECT  18.680 1.410 18.870 1.650 ;
        RECT  18.680 -0.400 21.720 0.400 ;
        RECT  21.720 -0.400 22.120 0.560 ;
        RECT  22.120 -0.400 23.180 0.400 ;
        RECT  23.180 -0.400 23.580 0.560 ;
        RECT  23.580 -0.400 24.420 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  23.250 2.170 23.650 2.570 ;
        RECT  22.940 2.250 23.250 2.490 ;
        RECT  22.700 1.260 22.940 4.010 ;
        RECT  22.540 1.260 22.700 1.660 ;
        RECT  22.500 3.610 22.700 4.010 ;
        RECT  21.570 3.690 22.500 3.930 ;
        RECT  21.720 2.240 22.430 2.640 ;
        RECT  21.480 1.270 21.720 2.640 ;
        RECT  21.360 2.920 21.570 3.930 ;
        RECT  20.890 1.270 21.480 1.510 ;
        RECT  20.890 2.400 21.480 2.640 ;
        RECT  21.170 2.920 21.360 4.370 ;
        RECT  19.960 1.880 21.200 2.120 ;
        RECT  21.120 3.690 21.170 4.370 ;
        RECT  14.520 4.130 21.120 4.370 ;
        RECT  20.730 1.110 20.890 1.510 ;
        RECT  20.650 2.400 20.890 3.240 ;
        RECT  20.490 0.670 20.730 1.510 ;
        RECT  20.550 3.000 20.650 3.240 ;
        RECT  20.390 3.000 20.550 3.400 ;
        RECT  18.970 0.670 20.490 0.910 ;
        RECT  20.150 3.000 20.390 3.850 ;
        RECT  18.630 3.610 20.150 3.850 ;
        RECT  19.440 1.200 20.130 1.440 ;
        RECT  19.720 1.880 19.960 2.730 ;
        RECT  19.440 3.080 19.790 3.320 ;
        RECT  19.200 1.200 19.440 3.320 ;
        RECT  18.110 1.970 19.200 2.210 ;
        RECT  18.310 2.500 18.830 2.740 ;
        RECT  18.070 2.500 18.310 3.850 ;
        RECT  17.790 1.130 18.110 2.210 ;
        RECT  15.000 3.610 18.070 3.850 ;
        RECT  17.710 1.130 17.790 3.330 ;
        RECT  17.550 1.970 17.710 3.330 ;
        RECT  17.290 3.090 17.550 3.330 ;
        RECT  17.020 2.200 17.260 2.600 ;
        RECT  16.950 2.360 17.020 2.600 ;
        RECT  16.710 2.360 16.950 3.330 ;
        RECT  15.550 3.090 16.710 3.330 ;
        RECT  16.070 1.220 16.470 1.460 ;
        RECT  16.070 2.570 16.230 2.810 ;
        RECT  15.830 1.220 16.070 2.810 ;
        RECT  15.310 0.940 15.550 3.330 ;
        RECT  14.120 2.280 15.310 2.520 ;
        RECT  15.090 2.900 15.310 3.140 ;
        RECT  14.760 3.420 15.000 3.850 ;
        RECT  14.720 1.330 14.960 1.980 ;
        RECT  12.950 3.420 14.760 3.660 ;
        RECT  13.470 1.330 14.720 1.570 ;
        RECT  14.280 3.940 14.520 4.370 ;
        RECT  12.430 3.940 14.280 4.180 ;
        RECT  13.880 1.850 14.120 2.520 ;
        RECT  13.230 1.020 13.470 3.130 ;
        RECT  12.750 1.020 13.230 1.260 ;
        RECT  12.760 2.840 12.950 3.660 ;
        RECT  12.710 1.600 12.760 3.660 ;
        RECT  12.520 1.600 12.710 3.080 ;
        RECT  12.380 1.600 12.520 1.840 ;
        RECT  10.770 2.840 12.520 3.080 ;
        RECT  12.190 3.470 12.430 4.180 ;
        RECT  12.140 1.100 12.380 1.840 ;
        RECT  10.350 3.470 12.190 3.710 ;
        RECT  11.210 1.100 12.140 1.340 ;
        RECT  10.810 0.940 11.210 1.340 ;
        RECT  8.980 4.120 10.970 4.360 ;
        RECT  10.230 0.910 10.470 1.310 ;
        RECT  10.230 3.310 10.350 3.710 ;
        RECT  9.990 0.910 10.230 3.710 ;
        RECT  9.470 0.910 9.710 3.830 ;
        RECT  9.270 0.910 9.470 1.310 ;
        RECT  9.270 3.360 9.470 3.830 ;
        RECT  6.750 3.360 9.270 3.600 ;
        RECT  8.990 2.190 9.190 3.080 ;
        RECT  8.750 0.750 8.990 3.080 ;
        RECT  8.740 3.880 8.980 4.360 ;
        RECT  8.450 0.750 8.750 1.100 ;
        RECT  8.740 2.440 8.750 2.880 ;
        RECT  3.010 3.880 8.740 4.120 ;
        RECT  8.230 2.420 8.470 2.820 ;
        RECT  7.180 0.860 8.450 1.100 ;
        RECT  7.530 2.580 8.230 2.820 ;
        RECT  7.330 2.580 7.530 3.080 ;
        RECT  7.150 2.350 7.330 3.080 ;
        RECT  7.150 1.380 7.310 1.620 ;
        RECT  6.940 0.670 7.180 1.100 ;
        RECT  7.090 1.380 7.150 3.080 ;
        RECT  6.910 1.380 7.090 2.590 ;
        RECT  5.900 0.670 6.940 0.910 ;
        RECT  6.790 2.190 6.910 2.590 ;
        RECT  6.510 3.040 6.750 3.600 ;
        RECT  6.510 1.230 6.570 1.470 ;
        RECT  6.270 1.230 6.510 3.600 ;
        RECT  6.170 1.230 6.270 1.470 ;
        RECT  3.770 3.360 6.270 3.600 ;
        RECT  5.890 2.840 5.990 3.080 ;
        RECT  5.650 1.230 5.890 3.080 ;
        RECT  5.290 1.230 5.650 1.470 ;
        RECT  5.590 2.840 5.650 3.080 ;
        RECT  4.290 2.830 4.510 3.070 ;
        RECT  4.050 1.390 4.290 3.070 ;
        RECT  3.810 1.390 4.050 2.540 ;
        RECT  3.530 3.180 3.770 3.600 ;
        RECT  3.530 0.680 3.690 0.920 ;
        RECT  3.290 0.680 3.530 3.600 ;
        RECT  2.770 1.330 3.010 4.120 ;
        RECT  2.710 1.330 2.770 1.740 ;
        RECT  2.610 2.990 2.770 3.390 ;
        RECT  1.960 3.670 2.360 4.260 ;
        RECT  2.030 1.340 2.130 1.740 ;
        RECT  2.030 2.980 2.110 3.380 ;
        RECT  1.790 1.340 2.030 3.380 ;
        RECT  0.570 3.670 1.960 3.910 ;
        RECT  1.730 1.340 1.790 1.740 ;
        RECT  1.710 2.980 1.790 3.380 ;
        RECT  0.400 1.340 0.570 1.740 ;
        RECT  0.400 2.980 0.570 3.910 ;
        RECT  0.330 1.340 0.400 3.910 ;
        RECT  0.160 1.340 0.330 3.390 ;
    END
END SEDFFHQX2

MACRO SEDFFHQX1
    CLASS CORE ;
    FOREIGN SEDFFHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SEDFFHQXL ;
    SIZE 23.100 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.530 0.720 2.180 1.040 ;
        RECT  2.180 0.710 2.440 1.040 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.710 2.010 0.860 2.640 ;
        RECT  0.860 2.010 1.120 2.650 ;
        RECT  1.120 2.010 1.160 2.640 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.980 1.260 22.530 1.540 ;
        RECT  22.530 1.260 22.650 1.700 ;
        RECT  22.530 3.060 22.690 3.460 ;
        RECT  22.650 1.260 22.690 1.840 ;
        RECT  22.690 1.260 22.930 3.460 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.590 1.420 8.120 1.660 ;
        RECT  8.120 1.270 8.370 1.660 ;
        RECT  8.370 1.270 8.380 1.530 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.820 1.830 5.120 2.090 ;
        RECT  5.120 1.730 5.520 2.130 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  11.390 1.740 11.910 2.140 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.960 5.440 ;
        RECT  0.960 4.480 1.360 5.440 ;
        RECT  1.360 4.640 5.020 5.440 ;
        RECT  5.020 4.480 5.420 5.440 ;
        RECT  5.420 4.640 7.940 5.440 ;
        RECT  7.940 4.480 8.340 5.440 ;
        RECT  8.340 4.640 11.820 5.440 ;
        RECT  11.820 3.840 12.220 5.440 ;
        RECT  12.220 4.640 14.710 5.440 ;
        RECT  14.710 4.480 15.110 5.440 ;
        RECT  15.110 4.640 20.190 5.440 ;
        RECT  20.190 4.590 20.200 5.440 ;
        RECT  20.200 4.480 20.600 5.440 ;
        RECT  20.600 4.590 21.770 5.440 ;
        RECT  21.770 4.480 22.170 5.440 ;
        RECT  22.170 4.590 22.180 5.440 ;
        RECT  22.180 4.640 23.100 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 4.640 0.400 ;
        RECT  4.640 -0.400 5.040 0.560 ;
        RECT  5.040 -0.400 8.000 0.400 ;
        RECT  8.000 -0.400 8.010 0.870 ;
        RECT  8.010 -0.400 8.410 0.990 ;
        RECT  8.410 -0.400 8.420 0.870 ;
        RECT  8.420 -0.400 11.980 0.400 ;
        RECT  11.980 -0.400 12.380 0.560 ;
        RECT  12.380 -0.400 14.650 0.400 ;
        RECT  14.650 -0.400 15.050 0.910 ;
        RECT  15.050 -0.400 17.360 0.400 ;
        RECT  17.360 -0.400 17.600 1.320 ;
        RECT  17.600 -0.400 20.350 0.400 ;
        RECT  20.350 -0.400 20.590 1.190 ;
        RECT  20.590 -0.400 21.770 0.400 ;
        RECT  21.770 -0.400 22.170 0.560 ;
        RECT  22.170 -0.400 23.100 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  22.010 2.260 22.410 2.660 ;
        RECT  21.490 2.340 22.010 2.580 ;
        RECT  21.430 1.040 21.490 3.640 ;
        RECT  21.250 1.040 21.430 4.300 ;
        RECT  21.030 1.040 21.250 1.440 ;
        RECT  21.030 3.400 21.250 4.300 ;
        RECT  20.360 3.400 21.030 3.640 ;
        RECT  20.070 2.030 20.920 2.430 ;
        RECT  19.960 2.920 20.360 3.640 ;
        RECT  19.830 0.670 20.070 2.610 ;
        RECT  19.920 3.400 19.960 3.640 ;
        RECT  19.680 3.400 19.920 4.370 ;
        RECT  18.820 0.670 19.830 0.910 ;
        RECT  19.260 2.370 19.830 2.610 ;
        RECT  15.630 4.130 19.680 4.370 ;
        RECT  19.380 1.250 19.540 1.490 ;
        RECT  19.140 1.250 19.380 2.120 ;
        RECT  19.020 2.370 19.260 3.430 ;
        RECT  18.740 1.880 19.140 2.120 ;
        RECT  18.500 1.880 18.740 3.850 ;
        RECT  18.400 2.340 18.500 2.740 ;
        RECT  16.160 3.610 18.500 3.850 ;
        RECT  18.120 1.130 18.460 1.530 ;
        RECT  18.120 3.090 18.220 3.330 ;
        RECT  17.880 1.130 18.120 3.330 ;
        RECT  17.820 3.090 17.880 3.330 ;
        RECT  17.300 1.960 17.540 3.140 ;
        RECT  15.860 2.900 17.300 3.140 ;
        RECT  16.400 0.820 16.800 1.220 ;
        RECT  16.380 2.380 16.580 2.620 ;
        RECT  16.380 0.980 16.400 1.220 ;
        RECT  16.140 0.980 16.380 2.620 ;
        RECT  15.920 3.420 16.160 3.850 ;
        RECT  13.240 3.420 15.920 3.660 ;
        RECT  15.620 0.920 15.860 3.140 ;
        RECT  15.390 3.940 15.630 4.370 ;
        RECT  14.890 2.900 15.620 3.140 ;
        RECT  12.720 3.940 15.390 4.180 ;
        RECT  15.050 1.150 15.290 1.820 ;
        RECT  13.920 1.150 15.050 1.390 ;
        RECT  14.880 2.320 14.890 3.140 ;
        RECT  14.650 2.240 14.880 3.140 ;
        RECT  14.480 2.240 14.650 2.640 ;
        RECT  13.680 0.930 13.920 3.140 ;
        RECT  13.310 0.930 13.680 1.170 ;
        RECT  13.530 2.740 13.680 3.140 ;
        RECT  13.240 1.510 13.400 1.750 ;
        RECT  13.000 1.510 13.240 3.660 ;
        RECT  12.660 1.510 13.000 1.750 ;
        RECT  11.000 2.840 13.000 3.080 ;
        RECT  12.480 3.360 12.720 4.180 ;
        RECT  12.420 1.220 12.660 1.750 ;
        RECT  10.610 3.360 12.480 3.600 ;
        RECT  11.770 1.220 12.420 1.460 ;
        RECT  11.370 1.060 11.770 1.460 ;
        RECT  10.800 3.880 11.200 4.280 ;
        RECT  10.610 0.910 10.910 1.310 ;
        RECT  3.030 3.880 10.800 4.120 ;
        RECT  10.370 0.910 10.610 3.600 ;
        RECT  10.210 2.980 10.370 3.380 ;
        RECT  9.890 0.910 10.030 1.310 ;
        RECT  9.770 0.910 9.890 3.100 ;
        RECT  9.650 0.910 9.770 3.600 ;
        RECT  9.630 0.910 9.650 1.310 ;
        RECT  9.530 2.780 9.650 3.600 ;
        RECT  6.810 3.360 9.530 3.600 ;
        RECT  9.190 1.920 9.350 2.320 ;
        RECT  9.190 0.770 9.290 1.170 ;
        RECT  8.950 0.770 9.190 3.110 ;
        RECT  8.890 0.770 8.950 1.170 ;
        RECT  8.710 2.870 8.950 3.110 ;
        RECT  8.250 2.060 8.650 2.460 ;
        RECT  7.550 2.220 8.250 2.460 ;
        RECT  7.310 2.220 7.550 3.110 ;
        RECT  7.310 0.670 7.530 1.070 ;
        RECT  7.150 0.670 7.310 3.110 ;
        RECT  7.070 0.670 7.150 2.460 ;
        RECT  6.830 2.030 7.070 2.460 ;
        RECT  6.550 2.960 6.810 3.600 ;
        RECT  6.550 1.040 6.790 1.440 ;
        RECT  6.310 1.040 6.550 3.600 ;
        RECT  3.810 3.360 6.310 3.600 ;
        RECT  5.790 1.030 6.030 3.080 ;
        RECT  5.590 1.030 5.790 1.440 ;
        RECT  5.630 2.840 5.790 3.080 ;
        RECT  5.510 1.040 5.590 1.440 ;
        RECT  4.330 2.830 4.550 3.070 ;
        RECT  4.330 1.340 4.360 1.740 ;
        RECT  4.090 1.340 4.330 3.070 ;
        RECT  3.960 1.340 4.090 1.740 ;
        RECT  3.910 2.150 4.090 2.660 ;
        RECT  3.630 3.050 3.810 3.600 ;
        RECT  3.630 0.680 3.650 0.920 ;
        RECT  3.390 0.680 3.630 3.600 ;
        RECT  3.250 0.680 3.390 0.920 ;
        RECT  2.950 2.990 3.030 4.120 ;
        RECT  2.950 1.340 2.990 1.740 ;
        RECT  2.790 1.340 2.950 4.120 ;
        RECT  2.710 1.340 2.790 3.390 ;
        RECT  2.590 1.340 2.710 1.740 ;
        RECT  2.630 2.990 2.710 3.390 ;
        RECT  2.000 3.670 2.400 4.250 ;
        RECT  2.050 2.980 2.130 3.380 ;
        RECT  2.050 1.340 2.110 1.740 ;
        RECT  1.810 1.340 2.050 3.380 ;
        RECT  0.570 3.670 2.000 3.910 ;
        RECT  1.710 1.340 1.810 1.740 ;
        RECT  1.730 2.980 1.810 3.380 ;
        RECT  0.400 1.340 0.570 1.740 ;
        RECT  0.400 2.980 0.570 3.910 ;
        RECT  0.330 1.340 0.400 3.910 ;
        RECT  0.160 1.340 0.330 3.390 ;
    END
END SEDFFHQX1

MACRO SEDFFXL
    CLASS CORE ;
    FOREIGN SEDFFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.390 2.240 3.850 2.660 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.390 1.600 2.650 ;
        RECT  1.600 2.250 2.000 2.650 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.840 1.400 18.020 1.830 ;
        RECT  17.910 2.620 18.030 3.240 ;
        RECT  18.020 1.400 18.030 2.090 ;
        RECT  18.030 1.400 18.270 3.240 ;
        RECT  18.270 1.830 18.280 2.090 ;
        RECT  18.270 2.620 18.310 3.240 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.450 3.510 16.720 3.990 ;
        RECT  16.720 3.500 16.850 3.990 ;
        RECT  16.850 3.500 16.960 3.770 ;
        RECT  16.570 0.740 16.970 1.110 ;
        RECT  16.960 3.500 17.280 3.740 ;
        RECT  16.970 0.870 17.280 1.110 ;
        RECT  17.280 0.870 17.520 3.740 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.470 3.750 0.770 4.150 ;
        RECT  0.770 3.510 1.010 4.150 ;
        RECT  1.010 3.510 1.120 3.770 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.400 2.250 4.800 2.630 ;
        RECT  4.800 2.390 4.820 2.630 ;
        RECT  4.820 2.390 5.080 2.650 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  10.010 1.830 10.520 2.230 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.300 5.440 ;
        RECT  1.300 4.050 1.700 5.440 ;
        RECT  1.700 4.640 2.920 5.440 ;
        RECT  2.920 4.130 3.320 5.440 ;
        RECT  3.320 4.640 9.340 5.440 ;
        RECT  9.340 4.480 10.940 5.440 ;
        RECT  10.940 4.640 12.200 5.440 ;
        RECT  12.200 4.480 13.180 5.440 ;
        RECT  13.180 4.640 15.630 5.440 ;
        RECT  15.630 3.220 16.030 5.440 ;
        RECT  16.030 4.600 17.240 5.440 ;
        RECT  17.240 4.480 17.640 5.440 ;
        RECT  17.640 4.640 18.480 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.360 0.400 ;
        RECT  0.360 -0.400 0.760 0.560 ;
        RECT  0.760 -0.400 3.330 0.400 ;
        RECT  3.330 -0.400 3.730 0.850 ;
        RECT  3.730 -0.400 10.730 0.400 ;
        RECT  10.730 -0.400 11.150 1.020 ;
        RECT  11.150 -0.400 12.870 0.400 ;
        RECT  12.870 -0.400 12.880 0.830 ;
        RECT  12.880 -0.400 13.280 1.030 ;
        RECT  13.280 -0.400 13.290 0.830 ;
        RECT  13.290 -0.400 15.770 0.400 ;
        RECT  15.770 -0.400 16.010 1.620 ;
        RECT  16.010 -0.400 17.890 0.400 ;
        RECT  17.890 -0.400 18.290 0.560 ;
        RECT  18.290 -0.400 18.480 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.970 2.160 17.040 3.140 ;
        RECT  16.730 1.380 16.970 3.140 ;
        RECT  16.570 1.380 16.730 1.780 ;
        RECT  16.500 2.740 16.730 3.140 ;
        RECT  15.310 2.740 16.500 2.980 ;
        RECT  15.490 2.070 16.400 2.470 ;
        RECT  15.250 0.690 15.490 2.470 ;
        RECT  15.070 2.740 15.310 4.180 ;
        RECT  14.210 0.690 15.250 0.930 ;
        RECT  14.590 2.230 15.250 2.470 ;
        RECT  7.390 3.940 15.070 4.180 ;
        RECT  14.110 1.250 14.970 1.490 ;
        RECT  14.350 2.230 14.590 3.660 ;
        RECT  14.130 3.260 14.350 3.660 ;
        RECT  13.890 1.250 14.110 2.740 ;
        RECT  13.870 1.250 13.890 3.660 ;
        RECT  13.650 2.500 13.870 3.660 ;
        RECT  9.080 3.420 13.650 3.660 ;
        RECT  13.090 1.420 13.330 3.140 ;
        RECT  12.540 1.420 13.090 1.660 ;
        RECT  12.300 2.900 13.090 3.140 ;
        RECT  11.840 2.330 12.810 2.570 ;
        RECT  12.400 1.260 12.540 1.660 ;
        RECT  12.140 0.670 12.400 1.660 ;
        RECT  12.000 0.670 12.140 0.910 ;
        RECT  11.710 2.330 11.840 3.070 ;
        RECT  11.470 1.240 11.710 3.070 ;
        RECT  9.600 2.830 11.470 3.070 ;
        RECT  10.990 1.310 11.230 2.290 ;
        RECT  10.460 1.310 10.990 1.550 ;
        RECT  10.220 0.670 10.460 1.550 ;
        RECT  8.490 0.670 10.220 0.910 ;
        RECT  9.080 1.320 9.940 1.560 ;
        RECT  9.360 2.150 9.600 3.070 ;
        RECT  8.840 1.320 9.080 3.660 ;
        RECT  7.380 1.710 8.840 1.950 ;
        RECT  8.320 3.420 8.840 3.660 ;
        RECT  8.250 0.670 8.490 1.090 ;
        RECT  8.250 2.730 8.410 3.130 ;
        RECT  8.080 0.850 8.250 1.090 ;
        RECT  8.010 2.230 8.250 3.130 ;
        RECT  7.680 0.850 8.080 1.430 ;
        RECT  7.100 2.230 8.010 2.470 ;
        RECT  7.100 1.190 7.680 1.430 ;
        RECT  7.130 2.800 7.530 3.200 ;
        RECT  7.150 3.480 7.390 4.180 ;
        RECT  4.300 0.680 7.200 0.920 ;
        RECT  6.990 3.480 7.150 3.880 ;
        RECT  6.710 2.960 7.130 3.200 ;
        RECT  6.860 1.190 7.100 2.470 ;
        RECT  6.470 2.960 6.710 4.260 ;
        RECT  4.370 4.020 6.470 4.260 ;
        RECT  3.750 3.500 6.190 3.740 ;
        RECT  6.020 1.730 6.180 2.010 ;
        RECT  5.780 1.730 6.020 3.170 ;
        RECT  3.090 1.200 5.860 1.440 ;
        RECT  2.610 1.730 5.780 1.970 ;
        RECT  5.390 2.930 5.780 3.170 ;
        RECT  3.080 2.970 4.340 3.210 ;
        RECT  3.510 3.500 3.750 3.850 ;
        RECT  2.570 3.610 3.510 3.850 ;
        RECT  2.850 0.690 3.090 1.440 ;
        RECT  2.760 2.250 3.080 3.210 ;
        RECT  2.310 0.690 2.850 0.930 ;
        RECT  2.680 2.250 2.760 2.490 ;
        RECT  2.570 2.970 2.760 3.210 ;
        RECT  2.370 1.210 2.610 1.970 ;
        RECT  2.170 2.970 2.570 3.320 ;
        RECT  2.170 3.610 2.570 4.140 ;
        RECT  0.570 1.210 2.370 1.450 ;
        RECT  1.190 2.970 2.170 3.210 ;
        RECT  1.190 1.730 2.130 1.970 ;
        RECT  0.950 1.730 1.190 3.210 ;
        RECT  0.490 1.210 0.570 1.800 ;
        RECT  0.250 1.210 0.490 3.380 ;
        RECT  0.170 1.400 0.250 1.800 ;
    END
END SEDFFXL

MACRO SEDFFX4
    CLASS CORE ;
    FOREIGN SEDFFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SEDFFXL ;
    SIZE 23.760 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 2.390 3.760 2.650 ;
        RECT  3.760 2.390 3.790 2.630 ;
        RECT  3.790 2.240 4.190 2.630 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.390 1.600 2.650 ;
        RECT  1.600 2.250 2.000 2.650 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  22.550 1.250 22.570 2.660 ;
        RECT  22.570 1.250 22.970 3.270 ;
        RECT  22.970 1.250 22.990 2.660 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.030 2.260 21.230 3.270 ;
        RECT  21.230 1.250 21.430 3.270 ;
        RECT  21.430 1.250 21.670 2.660 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.470 3.750 0.770 4.150 ;
        RECT  0.770 3.510 1.010 4.150 ;
        RECT  1.010 3.510 1.120 3.770 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.230 2.930 5.390 3.170 ;
        RECT  5.390 2.400 5.480 3.170 ;
        RECT  5.480 2.390 5.630 3.170 ;
        RECT  5.630 2.390 5.740 2.650 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  10.320 1.830 11.020 2.230 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.480 5.440 ;
        RECT  1.480 3.780 1.880 5.440 ;
        RECT  1.880 4.640 3.480 5.440 ;
        RECT  3.480 4.020 3.880 5.440 ;
        RECT  3.880 4.640 9.580 5.440 ;
        RECT  9.580 4.480 9.980 5.440 ;
        RECT  9.980 4.640 11.140 5.440 ;
        RECT  11.140 4.480 11.540 5.440 ;
        RECT  11.540 4.640 13.640 5.440 ;
        RECT  13.640 4.480 14.040 5.440 ;
        RECT  14.040 4.640 16.390 5.440 ;
        RECT  16.390 4.480 16.790 5.440 ;
        RECT  16.790 4.640 18.790 5.440 ;
        RECT  18.790 4.480 19.190 5.440 ;
        RECT  19.190 4.640 20.360 5.440 ;
        RECT  20.360 4.120 20.760 5.440 ;
        RECT  20.760 4.640 21.800 5.440 ;
        RECT  21.800 4.130 22.200 5.440 ;
        RECT  22.200 4.640 23.190 5.440 ;
        RECT  23.190 4.160 23.590 5.440 ;
        RECT  23.590 4.640 23.760 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.360 0.400 ;
        RECT  0.360 -0.400 0.760 0.560 ;
        RECT  0.760 -0.400 3.450 0.400 ;
        RECT  3.450 -0.400 3.850 0.920 ;
        RECT  3.850 -0.400 11.210 0.400 ;
        RECT  11.210 -0.400 11.450 1.030 ;
        RECT  11.450 -0.400 13.870 0.400 ;
        RECT  13.870 -0.400 14.270 1.040 ;
        RECT  14.270 -0.400 16.340 0.400 ;
        RECT  16.340 -0.400 16.740 0.560 ;
        RECT  16.740 -0.400 19.100 0.400 ;
        RECT  19.100 -0.400 19.500 1.610 ;
        RECT  19.500 -0.400 20.600 0.400 ;
        RECT  20.600 -0.400 21.000 0.960 ;
        RECT  21.000 -0.400 21.910 0.400 ;
        RECT  21.910 -0.400 22.310 0.970 ;
        RECT  22.310 -0.400 23.200 0.400 ;
        RECT  23.200 -0.400 23.600 0.970 ;
        RECT  23.600 -0.400 23.760 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  23.230 2.190 23.470 3.840 ;
        RECT  19.940 3.600 23.230 3.840 ;
        RECT  20.220 1.460 20.460 2.960 ;
        RECT  19.820 0.800 20.220 1.700 ;
        RECT  19.940 2.720 20.220 2.960 ;
        RECT  18.800 1.940 19.980 2.340 ;
        RECT  19.540 2.720 19.940 4.120 ;
        RECT  19.280 2.720 19.540 2.960 ;
        RECT  19.040 2.670 19.280 4.180 ;
        RECT  16.030 3.940 19.040 4.180 ;
        RECT  18.560 0.940 18.800 3.660 ;
        RECT  18.010 0.940 18.560 1.180 ;
        RECT  15.460 3.420 18.560 3.660 ;
        RECT  18.080 1.500 18.320 2.860 ;
        RECT  17.810 2.620 18.080 2.860 ;
        RECT  17.610 0.780 18.010 1.180 ;
        RECT  17.410 2.620 17.810 3.060 ;
        RECT  14.500 1.580 17.720 1.820 ;
        RECT  15.470 0.940 17.610 1.180 ;
        RECT  15.060 2.620 17.410 2.860 ;
        RECT  15.790 3.940 16.030 4.370 ;
        RECT  14.890 4.130 15.790 4.370 ;
        RECT  15.070 0.780 15.470 1.180 ;
        RECT  15.220 3.420 15.460 3.850 ;
        RECT  14.980 2.620 15.060 3.070 ;
        RECT  14.740 2.620 14.980 3.660 ;
        RECT  14.650 3.940 14.890 4.370 ;
        RECT  9.310 3.420 14.740 3.660 ;
        RECT  7.740 3.940 14.650 4.180 ;
        RECT  14.260 1.340 14.500 3.140 ;
        RECT  13.040 1.340 14.260 1.580 ;
        RECT  13.120 2.900 14.260 3.140 ;
        RECT  13.740 2.170 13.980 2.580 ;
        RECT  12.350 2.170 13.740 2.410 ;
        RECT  12.700 2.830 13.120 3.140 ;
        RECT  12.880 1.180 13.040 1.580 ;
        RECT  12.640 0.680 12.880 1.580 ;
        RECT  12.250 0.680 12.640 0.920 ;
        RECT  12.240 2.170 12.350 3.060 ;
        RECT  12.000 1.380 12.240 3.060 ;
        RECT  9.830 2.820 12.000 3.060 ;
        RECT  11.510 1.310 11.750 2.350 ;
        RECT  10.970 1.310 11.510 1.550 ;
        RECT  10.730 0.670 10.970 1.550 ;
        RECT  9.140 0.670 10.730 0.910 ;
        RECT  9.840 1.300 10.490 1.540 ;
        RECT  9.600 1.300 9.840 1.960 ;
        RECT  9.590 2.210 9.830 3.060 ;
        RECT  9.310 1.720 9.600 1.960 ;
        RECT  9.070 1.720 9.310 3.660 ;
        RECT  8.900 0.670 9.140 1.120 ;
        RECT  7.780 1.720 9.070 1.960 ;
        RECT  8.700 3.420 9.070 3.660 ;
        RECT  8.570 0.880 8.900 1.120 ;
        RECT  8.530 2.860 8.790 3.100 ;
        RECT  8.170 0.880 8.570 1.440 ;
        RECT  8.290 2.250 8.530 3.100 ;
        RECT  7.500 2.250 8.290 2.490 ;
        RECT  7.500 1.200 8.170 1.440 ;
        RECT  7.580 2.770 7.980 3.170 ;
        RECT  4.790 0.680 7.750 0.920 ;
        RECT  7.500 3.680 7.740 4.180 ;
        RECT  7.220 2.930 7.580 3.170 ;
        RECT  7.260 1.200 7.500 2.490 ;
        RECT  6.980 2.930 7.220 4.260 ;
        RECT  4.930 4.020 6.980 4.260 ;
        RECT  6.500 1.720 6.720 2.010 ;
        RECT  3.100 3.500 6.700 3.740 ;
        RECT  6.260 1.720 6.500 3.170 ;
        RECT  3.170 1.200 6.470 1.440 ;
        RECT  2.650 1.720 6.260 1.960 ;
        RECT  5.950 2.930 6.260 3.170 ;
        RECT  4.580 2.790 4.820 3.210 ;
        RECT  3.140 2.970 4.580 3.210 ;
        RECT  2.930 0.690 3.170 1.440 ;
        RECT  2.900 2.240 3.140 3.210 ;
        RECT  2.860 3.500 3.100 4.140 ;
        RECT  2.570 0.690 2.930 0.930 ;
        RECT  2.190 2.970 2.900 3.210 ;
        RECT  2.600 3.740 2.860 4.140 ;
        RECT  2.410 1.210 2.650 1.960 ;
        RECT  0.570 1.210 2.410 1.450 ;
        RECT  1.790 2.970 2.190 3.400 ;
        RECT  1.190 1.730 2.130 1.970 ;
        RECT  1.190 2.970 1.790 3.210 ;
        RECT  0.950 1.730 1.190 3.210 ;
        RECT  0.490 1.210 0.570 1.800 ;
        RECT  0.250 1.210 0.490 3.380 ;
        RECT  0.170 1.400 0.250 1.800 ;
    END
END SEDFFX4

MACRO SEDFFX2
    CLASS CORE ;
    FOREIGN SEDFFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SEDFFXL ;
    SIZE 20.460 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 2.390 3.520 2.650 ;
        RECT  3.520 2.240 3.980 2.660 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.290 2.250 1.690 2.650 ;
        RECT  1.690 2.390 1.780 2.650 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  19.890 1.250 19.910 1.650 ;
        RECT  19.890 3.070 20.010 4.050 ;
        RECT  19.910 1.250 20.010 1.820 ;
        RECT  20.010 1.250 20.250 4.050 ;
        RECT  20.250 3.070 20.290 4.050 ;
        RECT  20.250 1.250 20.290 1.960 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.460 2.820 18.590 3.230 ;
        RECT  18.590 2.660 18.690 3.230 ;
        RECT  18.630 1.260 18.690 1.820 ;
        RECT  18.690 1.260 18.930 3.230 ;
        RECT  18.930 1.260 19.030 1.820 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.470 3.750 0.770 4.150 ;
        RECT  0.770 3.520 0.860 4.150 ;
        RECT  0.860 3.510 1.010 4.150 ;
        RECT  1.010 3.510 1.120 3.770 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.400 2.250 4.820 2.490 ;
        RECT  4.820 2.250 5.080 2.650 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  10.050 1.940 10.100 2.340 ;
        RECT  10.100 1.830 10.360 2.340 ;
        RECT  10.360 1.940 10.450 2.340 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.480 5.440 ;
        RECT  1.480 3.780 1.880 5.440 ;
        RECT  1.880 4.640 3.110 5.440 ;
        RECT  3.110 4.020 3.510 5.440 ;
        RECT  3.510 4.640 9.280 5.440 ;
        RECT  9.280 4.480 10.880 5.440 ;
        RECT  10.880 4.640 12.180 5.440 ;
        RECT  12.180 4.480 13.240 5.440 ;
        RECT  13.240 4.640 15.700 5.440 ;
        RECT  15.700 4.480 17.240 5.440 ;
        RECT  17.240 4.600 19.130 5.440 ;
        RECT  19.130 4.130 19.530 5.440 ;
        RECT  19.530 4.640 20.460 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.360 0.400 ;
        RECT  0.360 -0.400 0.760 0.560 ;
        RECT  0.760 -0.400 3.440 0.400 ;
        RECT  3.440 -0.400 3.450 0.730 ;
        RECT  3.450 -0.400 3.850 0.850 ;
        RECT  3.850 -0.400 3.860 0.730 ;
        RECT  3.860 -0.400 10.730 0.400 ;
        RECT  10.730 -0.400 11.150 0.930 ;
        RECT  11.150 -0.400 12.730 0.400 ;
        RECT  12.730 -0.400 12.740 0.670 ;
        RECT  12.740 -0.400 13.140 0.870 ;
        RECT  13.140 -0.400 13.150 0.670 ;
        RECT  13.150 -0.400 15.300 0.400 ;
        RECT  15.300 -0.400 15.310 0.850 ;
        RECT  15.310 -0.400 15.710 1.050 ;
        RECT  15.710 -0.400 15.720 0.850 ;
        RECT  15.720 -0.400 17.240 0.400 ;
        RECT  17.240 -0.400 17.660 1.430 ;
        RECT  17.660 -0.400 19.240 0.400 ;
        RECT  19.240 -0.400 19.250 0.770 ;
        RECT  19.250 -0.400 19.650 0.970 ;
        RECT  19.650 -0.400 19.660 0.770 ;
        RECT  19.660 -0.400 20.460 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  19.400 2.250 19.640 3.850 ;
        RECT  18.160 3.610 19.400 3.850 ;
        RECT  18.160 1.140 18.210 2.530 ;
        RECT  17.970 1.140 18.160 3.980 ;
        RECT  17.920 2.290 17.970 3.980 ;
        RECT  17.630 3.580 17.920 3.980 ;
        RECT  16.970 1.820 17.640 2.220 ;
        RECT  16.880 3.740 17.630 3.980 ;
        RECT  16.730 1.550 16.970 2.990 ;
        RECT  16.480 3.740 16.880 4.180 ;
        RECT  16.230 1.550 16.730 1.790 ;
        RECT  16.410 2.750 16.730 2.990 ;
        RECT  16.080 2.060 16.480 2.460 ;
        RECT  7.260 3.940 16.480 4.180 ;
        RECT  16.120 2.750 16.410 3.150 ;
        RECT  15.830 1.340 16.230 1.790 ;
        RECT  15.880 2.750 16.120 3.580 ;
        RECT  15.350 2.220 16.080 2.460 ;
        RECT  14.510 3.340 15.880 3.580 ;
        RECT  14.420 1.340 15.830 1.580 ;
        RECT  15.110 2.220 15.350 2.740 ;
        RECT  14.250 2.500 15.110 2.740 ;
        RECT  13.210 1.860 14.660 2.100 ;
        RECT  14.110 3.260 14.510 3.660 ;
        RECT  14.020 1.100 14.420 1.580 ;
        RECT  13.850 2.500 14.250 2.900 ;
        RECT  13.610 2.500 13.850 3.660 ;
        RECT  8.820 3.420 13.610 3.660 ;
        RECT  12.970 1.410 13.210 3.140 ;
        RECT  12.430 1.410 12.970 1.660 ;
        RECT  12.190 2.900 12.970 3.140 ;
        RECT  11.720 2.330 12.690 2.570 ;
        RECT  12.270 1.260 12.430 1.660 ;
        RECT  12.030 0.670 12.270 1.660 ;
        RECT  11.480 0.670 12.030 0.910 ;
        RECT  11.610 2.330 11.720 3.080 ;
        RECT  11.370 1.380 11.610 3.080 ;
        RECT  9.340 2.840 11.370 3.080 ;
        RECT  10.850 1.310 11.090 2.340 ;
        RECT  10.460 1.310 10.850 1.550 ;
        RECT  10.220 0.670 10.460 1.550 ;
        RECT  8.480 0.670 10.220 0.910 ;
        RECT  9.510 1.310 9.940 1.550 ;
        RECT  9.270 1.310 9.510 1.870 ;
        RECT  9.100 2.150 9.340 3.080 ;
        RECT  8.820 1.630 9.270 1.870 ;
        RECT  8.580 1.630 8.820 3.660 ;
        RECT  7.320 1.720 8.580 1.960 ;
        RECT  8.220 3.420 8.580 3.660 ;
        RECT  8.240 0.670 8.480 1.110 ;
        RECT  8.140 2.840 8.300 3.080 ;
        RECT  8.080 0.870 8.240 1.110 ;
        RECT  7.900 2.250 8.140 3.080 ;
        RECT  7.680 0.870 8.080 1.440 ;
        RECT  7.040 2.250 7.900 2.490 ;
        RECT  7.040 1.200 7.680 1.440 ;
        RECT  7.100 2.760 7.500 3.160 ;
        RECT  7.020 3.480 7.260 4.180 ;
        RECT  4.710 0.680 7.200 0.920 ;
        RECT  6.740 2.920 7.100 3.160 ;
        RECT  6.800 1.200 7.040 2.490 ;
        RECT  6.500 2.920 6.740 4.260 ;
        RECT  4.450 4.020 6.500 4.260 ;
        RECT  2.730 3.500 6.220 3.740 ;
        RECT  6.020 1.730 6.180 2.010 ;
        RECT  5.780 1.730 6.020 3.170 ;
        RECT  3.170 1.200 5.860 1.440 ;
        RECT  2.650 1.730 5.780 1.970 ;
        RECT  5.470 2.930 5.780 3.170 ;
        RECT  4.310 0.670 4.710 0.920 ;
        RECT  3.130 2.970 4.530 3.210 ;
        RECT  2.930 0.690 3.170 1.440 ;
        RECT  2.890 2.280 3.130 3.210 ;
        RECT  2.310 0.690 2.930 0.930 ;
        RECT  2.190 2.970 2.890 3.210 ;
        RECT  2.490 3.500 2.730 4.140 ;
        RECT  2.410 1.210 2.650 1.970 ;
        RECT  2.230 3.740 2.490 4.140 ;
        RECT  0.570 1.210 2.410 1.450 ;
        RECT  1.790 2.970 2.190 3.400 ;
        RECT  1.050 1.730 2.140 1.970 ;
        RECT  1.050 2.970 1.790 3.210 ;
        RECT  0.810 1.730 1.050 3.210 ;
        RECT  0.490 1.210 0.570 1.800 ;
        RECT  0.250 1.210 0.490 3.380 ;
        RECT  0.170 1.400 0.250 1.800 ;
    END
END SEDFFX2

MACRO SEDFFX1
    CLASS CORE ;
    FOREIGN SEDFFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SEDFFXL ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.390 2.240 3.850 2.660 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.390 1.600 2.660 ;
        RECT  1.600 2.260 2.000 2.660 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.910 1.270 17.930 1.670 ;
        RECT  17.910 3.090 18.030 3.490 ;
        RECT  17.930 1.270 18.030 1.820 ;
        RECT  18.030 1.270 18.270 3.490 ;
        RECT  18.270 3.090 18.310 3.490 ;
        RECT  18.270 1.270 18.310 1.960 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.490 3.750 16.620 4.150 ;
        RECT  16.620 3.510 16.890 4.150 ;
        RECT  16.510 0.730 16.910 1.110 ;
        RECT  16.890 3.510 16.960 3.770 ;
        RECT  16.960 3.510 17.320 3.750 ;
        RECT  16.910 0.870 17.320 1.110 ;
        RECT  17.320 0.870 17.560 3.750 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.470 3.750 0.770 4.150 ;
        RECT  0.770 3.520 0.860 4.150 ;
        RECT  0.860 3.510 1.010 4.150 ;
        RECT  1.010 3.510 1.120 3.770 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.410 2.250 4.820 2.650 ;
        RECT  4.820 2.390 5.080 2.650 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  10.100 1.830 10.240 2.090 ;
        RECT  10.240 1.830 10.640 2.230 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.280 5.440 ;
        RECT  1.280 4.250 1.290 5.440 ;
        RECT  1.290 4.050 1.690 5.440 ;
        RECT  1.690 4.250 1.700 5.440 ;
        RECT  1.700 4.640 3.110 5.440 ;
        RECT  3.110 4.010 3.510 5.440 ;
        RECT  3.510 4.640 9.340 5.440 ;
        RECT  9.340 4.480 10.880 5.440 ;
        RECT  10.880 4.640 12.080 5.440 ;
        RECT  12.080 4.480 13.060 5.440 ;
        RECT  13.060 4.640 15.690 5.440 ;
        RECT  15.690 3.470 16.090 5.440 ;
        RECT  16.090 4.600 17.220 5.440 ;
        RECT  17.220 4.480 17.620 5.440 ;
        RECT  17.620 4.640 18.480 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.360 0.400 ;
        RECT  0.360 -0.400 0.760 0.560 ;
        RECT  0.760 -0.400 3.340 0.400 ;
        RECT  3.340 -0.400 3.740 0.940 ;
        RECT  3.740 -0.400 10.700 0.400 ;
        RECT  10.700 -0.400 10.940 1.000 ;
        RECT  10.940 -0.400 12.870 0.400 ;
        RECT  12.870 -0.400 12.880 0.830 ;
        RECT  12.880 -0.400 13.280 1.030 ;
        RECT  13.280 -0.400 13.290 0.830 ;
        RECT  13.290 -0.400 15.770 0.400 ;
        RECT  15.770 -0.400 16.010 1.480 ;
        RECT  16.010 -0.400 17.800 0.400 ;
        RECT  17.800 -0.400 18.200 0.560 ;
        RECT  18.200 -0.400 18.480 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.970 2.170 17.040 3.150 ;
        RECT  16.730 1.380 16.970 3.150 ;
        RECT  16.570 1.380 16.730 1.780 ;
        RECT  16.490 2.750 16.730 3.150 ;
        RECT  15.190 2.890 16.490 3.130 ;
        RECT  15.490 2.070 16.390 2.470 ;
        RECT  15.250 0.690 15.490 2.610 ;
        RECT  14.220 0.690 15.250 0.930 ;
        RECT  14.440 2.370 15.250 2.610 ;
        RECT  14.950 2.890 15.190 4.180 ;
        RECT  14.800 1.250 14.960 1.490 ;
        RECT  7.390 3.940 14.950 4.180 ;
        RECT  14.560 1.250 14.800 2.060 ;
        RECT  13.960 1.820 14.560 2.060 ;
        RECT  14.200 2.370 14.440 3.430 ;
        RECT  14.010 3.030 14.200 3.430 ;
        RECT  13.730 1.820 13.960 2.740 ;
        RECT  13.720 1.820 13.730 3.660 ;
        RECT  13.490 2.490 13.720 3.660 ;
        RECT  9.080 3.420 13.490 3.660 ;
        RECT  12.970 1.410 13.210 3.140 ;
        RECT  12.540 1.410 12.970 1.650 ;
        RECT  12.190 2.900 12.970 3.140 ;
        RECT  11.720 2.330 12.690 2.570 ;
        RECT  12.410 1.250 12.540 1.650 ;
        RECT  12.400 0.900 12.410 1.650 ;
        RECT  12.140 0.670 12.400 1.650 ;
        RECT  12.000 0.670 12.140 0.910 ;
        RECT  11.480 1.260 11.720 3.070 ;
        RECT  9.600 2.830 11.480 3.070 ;
        RECT  11.000 1.310 11.240 2.290 ;
        RECT  10.460 1.310 11.000 1.550 ;
        RECT  10.220 0.670 10.460 1.550 ;
        RECT  8.480 0.670 10.220 0.910 ;
        RECT  9.080 1.320 9.940 1.560 ;
        RECT  9.360 2.150 9.600 3.070 ;
        RECT  8.840 1.320 9.080 3.660 ;
        RECT  7.380 1.710 8.840 1.950 ;
        RECT  8.330 3.420 8.840 3.660 ;
        RECT  8.240 0.670 8.480 1.090 ;
        RECT  8.250 2.740 8.410 3.140 ;
        RECT  8.010 2.230 8.250 3.140 ;
        RECT  8.080 0.850 8.240 1.090 ;
        RECT  7.680 0.850 8.080 1.430 ;
        RECT  7.100 2.230 8.010 2.470 ;
        RECT  7.100 1.190 7.680 1.430 ;
        RECT  7.130 2.800 7.530 3.200 ;
        RECT  7.150 3.470 7.390 4.180 ;
        RECT  4.300 0.680 7.200 0.920 ;
        RECT  6.990 3.470 7.150 3.870 ;
        RECT  6.710 2.960 7.130 3.200 ;
        RECT  6.860 1.190 7.100 2.470 ;
        RECT  6.470 2.960 6.710 4.250 ;
        RECT  4.450 4.010 6.470 4.250 ;
        RECT  2.830 3.490 6.190 3.730 ;
        RECT  6.020 1.730 6.180 2.010 ;
        RECT  5.780 1.730 6.020 3.170 ;
        RECT  3.100 1.200 5.860 1.440 ;
        RECT  2.610 1.730 5.780 1.970 ;
        RECT  5.220 2.930 5.780 3.170 ;
        RECT  3.080 2.970 4.370 3.210 ;
        RECT  2.860 0.730 3.100 1.440 ;
        RECT  2.760 2.280 3.080 3.210 ;
        RECT  2.320 0.730 2.860 0.970 ;
        RECT  2.590 3.490 2.830 4.240 ;
        RECT  2.680 2.280 2.760 2.680 ;
        RECT  2.310 2.970 2.760 3.210 ;
        RECT  2.370 1.210 2.610 1.970 ;
        RECT  2.230 3.840 2.590 4.240 ;
        RECT  0.570 1.210 2.370 1.450 ;
        RECT  1.910 2.970 2.310 3.400 ;
        RECT  1.160 1.730 2.130 1.970 ;
        RECT  1.160 2.970 1.910 3.210 ;
        RECT  0.920 1.730 1.160 3.210 ;
        RECT  0.490 1.210 0.570 1.790 ;
        RECT  0.250 1.210 0.490 3.380 ;
        RECT  0.170 1.390 0.250 1.790 ;
    END
END SEDFFX1

MACRO SDFFTRXL
    CLASS CORE ;
    FOREIGN SDFFTRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.160 2.420 3.170 2.660 ;
        RECT  3.170 2.380 3.760 2.680 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.000 2.110 2.240 2.550 ;
        RECT  2.240 2.310 2.390 2.550 ;
        RECT  2.390 2.310 2.630 3.180 ;
        RECT  2.630 2.940 2.840 3.180 ;
        RECT  2.840 2.940 2.860 3.210 ;
        RECT  2.860 2.940 3.080 3.250 ;
        RECT  3.080 2.950 3.100 3.250 ;
        RECT  3.100 3.010 4.240 3.250 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.110 1.910 4.350 2.630 ;
        RECT  4.350 2.390 4.820 2.630 ;
        RECT  4.820 2.390 5.080 2.650 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.030 1.170 15.290 1.570 ;
        RECT  14.940 3.080 15.300 3.480 ;
        RECT  15.290 1.170 15.300 1.890 ;
        RECT  15.300 1.170 15.540 3.480 ;
        RECT  15.540 1.170 15.630 2.090 ;
        RECT  15.630 1.260 15.640 2.090 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.410 3.500 13.420 4.050 ;
        RECT  13.320 0.670 13.440 0.910 ;
        RECT  13.440 0.670 13.720 1.100 ;
        RECT  13.420 3.500 13.820 4.110 ;
        RECT  13.820 3.500 14.350 3.780 ;
        RECT  13.720 0.860 14.350 1.100 ;
        RECT  14.350 0.860 14.590 3.780 ;
        RECT  14.590 3.500 14.600 3.780 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.030 1.240 5.480 1.480 ;
        RECT  5.480 1.240 5.730 1.530 ;
        RECT  5.730 1.270 5.740 1.530 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.710 2.120 1.170 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.740 5.440 ;
        RECT  0.740 4.480 1.140 5.440 ;
        RECT  1.140 4.640 8.060 5.440 ;
        RECT  8.060 4.480 8.460 5.440 ;
        RECT  8.460 4.640 10.310 5.440 ;
        RECT  10.310 3.890 10.320 5.440 ;
        RECT  10.320 3.690 10.720 5.440 ;
        RECT  10.720 3.890 10.730 5.440 ;
        RECT  10.730 4.640 12.590 5.440 ;
        RECT  12.590 4.170 12.600 5.440 ;
        RECT  12.600 3.970 13.000 5.440 ;
        RECT  13.000 4.170 13.010 5.440 ;
        RECT  13.010 4.640 14.240 5.440 ;
        RECT  14.240 4.480 14.640 5.440 ;
        RECT  14.640 4.640 15.840 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        RECT  0.900 -0.400 1.300 0.560 ;
        RECT  1.300 -0.400 3.010 0.400 ;
        RECT  3.010 -0.400 3.410 0.560 ;
        RECT  3.410 -0.400 7.880 0.400 ;
        RECT  7.880 -0.400 7.890 0.730 ;
        RECT  7.890 -0.400 8.290 0.850 ;
        RECT  8.290 -0.400 8.300 0.730 ;
        RECT  8.300 -0.400 10.170 0.400 ;
        RECT  10.170 -0.400 10.410 1.150 ;
        RECT  10.410 -0.400 12.500 0.400 ;
        RECT  12.500 -0.400 12.900 0.560 ;
        RECT  12.900 -0.400 14.060 0.400 ;
        RECT  14.060 -0.400 14.460 0.560 ;
        RECT  14.460 -0.400 15.840 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  13.830 1.540 14.070 3.160 ;
        RECT  13.780 1.540 13.830 1.780 ;
        RECT  13.510 2.760 13.830 3.160 ;
        RECT  13.380 1.380 13.780 1.780 ;
        RECT  13.150 2.060 13.430 2.460 ;
        RECT  12.630 1.540 13.380 1.780 ;
        RECT  13.030 2.060 13.150 3.130 ;
        RECT  12.910 2.120 13.030 3.130 ;
        RECT  12.110 2.890 12.910 3.130 ;
        RECT  12.390 1.540 12.630 2.260 ;
        RECT  12.060 1.220 12.110 4.030 ;
        RECT  11.870 1.220 12.060 4.110 ;
        RECT  11.690 1.220 11.870 1.460 ;
        RECT  11.790 2.890 11.870 4.110 ;
        RECT  11.660 3.710 11.790 4.110 ;
        RECT  11.450 1.060 11.690 1.460 ;
        RECT  11.170 1.880 11.530 2.120 ;
        RECT  10.930 1.430 11.170 2.980 ;
        RECT  9.860 1.430 10.930 1.670 ;
        RECT  10.200 2.740 10.930 2.980 ;
        RECT  10.400 1.950 10.640 2.350 ;
        RECT  9.210 1.960 10.400 2.350 ;
        RECT  9.960 2.740 10.200 3.220 ;
        RECT  9.620 0.670 9.860 1.670 ;
        RECT  9.680 4.130 9.760 4.370 ;
        RECT  9.360 3.940 9.680 4.370 ;
        RECT  9.210 0.670 9.620 0.990 ;
        RECT  7.400 3.940 9.360 4.180 ;
        RECT  8.810 0.750 9.210 0.990 ;
        RECT  9.010 1.600 9.210 3.140 ;
        RECT  8.970 1.450 9.010 3.140 ;
        RECT  8.770 1.450 8.970 1.850 ;
        RECT  7.840 2.900 8.970 3.140 ;
        RECT  8.570 0.670 8.810 1.070 ;
        RECT  8.360 2.250 8.680 2.490 ;
        RECT  8.120 1.610 8.360 2.490 ;
        RECT  7.280 1.610 8.120 1.850 ;
        RECT  7.600 2.130 7.840 3.140 ;
        RECT  6.950 3.940 7.400 4.360 ;
        RECT  7.040 0.670 7.280 2.860 ;
        RECT  6.080 0.670 7.040 0.910 ;
        RECT  6.980 2.620 7.040 2.860 ;
        RECT  6.740 2.620 6.980 3.050 ;
        RECT  6.280 4.120 6.950 4.360 ;
        RECT  6.680 1.660 6.760 1.900 ;
        RECT  6.360 1.660 6.680 2.080 ;
        RECT  6.280 1.840 6.360 2.080 ;
        RECT  6.040 1.840 6.280 4.360 ;
        RECT  1.680 4.120 6.040 4.360 ;
        RECT  5.680 3.600 5.750 3.840 ;
        RECT  5.440 2.250 5.680 3.840 ;
        RECT  3.930 0.670 5.670 0.910 ;
        RECT  5.350 3.590 5.440 3.840 ;
        RECT  2.080 3.590 5.350 3.830 ;
        RECT  4.600 1.240 4.710 1.480 ;
        RECT  4.310 1.240 4.600 1.620 ;
        RECT  3.030 1.380 4.310 1.620 ;
        RECT  3.690 0.670 3.930 1.100 ;
        RECT  2.040 0.860 3.690 1.100 ;
        RECT  2.790 1.380 3.030 2.010 ;
        RECT  1.790 1.380 2.790 1.790 ;
        RECT  1.720 2.830 2.110 3.070 ;
        RECT  1.720 0.720 2.040 1.100 ;
        RECT  1.720 1.550 1.790 1.790 ;
        RECT  1.640 0.720 1.720 0.960 ;
        RECT  1.480 1.550 1.720 3.070 ;
        RECT  1.440 3.940 1.680 4.360 ;
        RECT  0.490 3.940 1.440 4.180 ;
        RECT  0.430 1.280 0.570 1.680 ;
        RECT  0.490 2.970 0.570 3.370 ;
        RECT  0.430 2.970 0.490 4.180 ;
        RECT  0.250 1.280 0.430 4.180 ;
        RECT  0.190 1.280 0.250 3.370 ;
        RECT  0.170 1.280 0.190 1.680 ;
        RECT  0.170 2.970 0.190 3.370 ;
    END
END SDFFTRXL

MACRO SDFFTRX4
    CLASS CORE ;
    FOREIGN SDFFTRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFTRXL ;
    SIZE 21.120 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.930 2.930 4.860 3.220 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.000 2.400 2.180 2.690 ;
        RECT  2.180 2.390 2.440 2.690 ;
        RECT  2.440 2.420 2.520 2.690 ;
        RECT  2.520 2.420 5.410 2.660 ;
        RECT  5.410 2.420 5.650 3.100 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.170 1.900 5.930 2.140 ;
        RECT  5.930 1.900 6.170 2.650 ;
        RECT  6.170 2.170 6.400 2.650 ;
        RECT  6.400 2.170 6.450 2.570 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  19.250 1.260 19.420 2.660 ;
        RECT  19.420 1.260 19.830 3.160 ;
        RECT  19.830 1.390 19.840 3.160 ;
        RECT  19.840 2.750 20.030 3.150 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.930 1.820 18.080 3.220 ;
        RECT  18.080 1.460 18.090 3.220 ;
        RECT  18.090 1.260 18.370 3.220 ;
        RECT  18.370 1.260 18.490 3.210 ;
        RECT  18.490 1.460 18.500 3.010 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.300 1.820 3.200 2.120 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.710 2.090 1.120 2.660 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.980 5.440 ;
        RECT  0.980 3.870 1.380 5.440 ;
        RECT  1.380 4.640 9.390 5.440 ;
        RECT  9.390 4.480 9.790 5.440 ;
        RECT  9.790 4.640 10.690 5.440 ;
        RECT  10.690 4.480 11.090 5.440 ;
        RECT  11.090 4.640 13.170 5.440 ;
        RECT  13.170 3.930 13.180 5.440 ;
        RECT  13.180 3.730 13.580 5.440 ;
        RECT  13.580 3.930 13.590 5.440 ;
        RECT  13.590 4.640 16.040 5.440 ;
        RECT  16.040 4.480 16.440 5.440 ;
        RECT  16.440 4.640 17.440 5.440 ;
        RECT  17.440 4.210 17.450 5.440 ;
        RECT  17.450 4.010 17.850 5.440 ;
        RECT  17.850 4.210 17.860 5.440 ;
        RECT  17.860 4.640 18.850 5.440 ;
        RECT  18.850 4.210 18.860 5.440 ;
        RECT  18.860 4.010 19.260 5.440 ;
        RECT  19.260 4.210 19.270 5.440 ;
        RECT  19.270 4.640 20.270 5.440 ;
        RECT  20.270 4.010 20.670 5.440 ;
        RECT  20.670 4.640 21.120 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        RECT  0.980 -0.400 1.380 0.560 ;
        RECT  1.380 -0.400 4.510 0.400 ;
        RECT  4.510 -0.400 4.910 0.560 ;
        RECT  4.910 -0.400 7.940 0.400 ;
        RECT  7.940 -0.400 7.950 1.240 ;
        RECT  7.950 -0.400 8.350 1.440 ;
        RECT  8.350 -0.400 8.360 1.240 ;
        RECT  8.360 -0.400 10.610 0.400 ;
        RECT  10.610 -0.400 10.620 1.110 ;
        RECT  10.620 -0.400 11.020 1.310 ;
        RECT  11.020 -0.400 11.030 1.110 ;
        RECT  11.030 -0.400 13.150 0.400 ;
        RECT  13.150 -0.400 13.160 1.130 ;
        RECT  13.160 -0.400 13.560 1.330 ;
        RECT  13.560 -0.400 13.570 1.130 ;
        RECT  13.570 -0.400 15.890 0.400 ;
        RECT  15.890 -0.400 16.290 0.560 ;
        RECT  16.290 -0.400 17.440 0.400 ;
        RECT  17.440 -0.400 17.450 0.780 ;
        RECT  17.450 -0.400 17.850 0.980 ;
        RECT  17.850 -0.400 17.860 0.780 ;
        RECT  17.860 -0.400 18.750 0.400 ;
        RECT  18.750 -0.400 18.760 0.780 ;
        RECT  18.760 -0.400 19.160 0.980 ;
        RECT  19.160 -0.400 19.170 0.780 ;
        RECT  19.170 -0.400 20.060 0.400 ;
        RECT  20.060 -0.400 20.070 0.780 ;
        RECT  20.070 -0.400 20.470 0.980 ;
        RECT  20.470 -0.400 20.480 0.780 ;
        RECT  20.480 -0.400 21.120 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  20.310 2.070 20.550 3.730 ;
        RECT  20.140 2.070 20.310 2.470 ;
        RECT  17.660 3.490 20.310 3.730 ;
        RECT  17.420 1.380 17.660 3.730 ;
        RECT  17.110 1.380 17.420 1.620 ;
        RECT  16.710 2.910 17.420 3.310 ;
        RECT  16.740 2.110 17.140 2.510 ;
        RECT  16.710 1.220 17.110 1.620 ;
        RECT  16.430 2.110 16.740 2.350 ;
        RECT  15.770 3.070 16.710 3.310 ;
        RECT  16.190 1.370 16.430 2.350 ;
        RECT  14.780 1.370 16.190 1.610 ;
        RECT  15.530 3.070 15.770 3.720 ;
        RECT  15.240 1.890 15.440 2.130 ;
        RECT  15.000 1.890 15.240 4.360 ;
        RECT  14.100 4.120 15.000 4.360 ;
        RECT  14.720 1.210 14.780 1.610 ;
        RECT  14.480 1.210 14.720 3.460 ;
        RECT  14.380 1.210 14.480 1.610 ;
        RECT  12.360 2.090 14.480 2.330 ;
        RECT  13.860 3.210 14.100 4.360 ;
        RECT  12.880 3.210 13.860 3.450 ;
        RECT  12.640 3.210 12.880 4.080 ;
        RECT  10.390 3.840 12.640 4.080 ;
        RECT  12.340 2.090 12.360 3.560 ;
        RECT  12.100 1.060 12.340 3.560 ;
        RECT  11.940 1.060 12.100 1.460 ;
        RECT  11.960 3.160 12.100 3.560 ;
        RECT  11.420 1.590 11.660 3.050 ;
        RECT  10.260 1.590 11.420 1.830 ;
        RECT  10.210 2.810 11.420 3.050 ;
        RECT  9.320 2.110 11.140 2.510 ;
        RECT  9.990 3.780 10.390 4.180 ;
        RECT  10.100 1.030 10.260 1.830 ;
        RECT  10.020 0.670 10.100 1.830 ;
        RECT  9.860 0.670 10.020 1.430 ;
        RECT  8.040 3.940 9.990 4.180 ;
        RECT  9.290 0.670 9.860 0.910 ;
        RECT  9.080 1.200 9.320 2.910 ;
        RECT  8.710 1.200 9.080 1.600 ;
        RECT  9.070 2.670 9.080 2.910 ;
        RECT  8.690 2.670 9.070 3.070 ;
        RECT  8.400 1.880 8.800 2.280 ;
        RECT  8.310 2.660 8.690 3.080 ;
        RECT  7.520 1.960 8.400 2.200 ;
        RECT  8.010 2.670 8.310 3.070 ;
        RECT  7.800 3.940 8.040 4.370 ;
        RECT  6.790 4.130 7.800 4.370 ;
        RECT  7.310 0.860 7.520 3.690 ;
        RECT  7.280 0.860 7.310 3.850 ;
        RECT  6.610 0.860 7.280 1.100 ;
        RECT  7.070 3.450 7.280 3.850 ;
        RECT  6.790 1.610 7.000 3.170 ;
        RECT  6.760 1.610 6.790 4.370 ;
        RECT  6.690 1.610 6.760 1.850 ;
        RECT  6.550 2.930 6.760 4.370 ;
        RECT  6.450 1.380 6.690 1.850 ;
        RECT  3.710 1.380 6.450 1.620 ;
        RECT  6.030 3.490 6.270 4.190 ;
        RECT  4.230 0.860 6.250 1.100 ;
        RECT  3.550 3.490 6.030 3.730 ;
        RECT  2.860 4.010 5.590 4.250 ;
        RECT  3.990 0.790 4.230 1.100 ;
        RECT  2.770 0.790 3.990 1.030 ;
        RECT  3.470 1.310 3.710 1.620 ;
        RECT  3.230 3.460 3.550 3.730 ;
        RECT  2.490 1.310 3.470 1.550 ;
        RECT  3.150 3.460 3.230 3.700 ;
        RECT  2.620 3.460 2.860 4.250 ;
        RECT  2.390 3.460 2.620 3.700 ;
        RECT  2.250 0.860 2.490 1.550 ;
        RECT  1.970 4.110 2.340 4.350 ;
        RECT  0.570 0.860 2.250 1.100 ;
        RECT  1.730 1.390 1.970 1.790 ;
        RECT  1.730 2.990 1.970 4.350 ;
        RECT  1.720 1.550 1.730 1.790 ;
        RECT  1.720 2.990 1.730 3.230 ;
        RECT  1.480 1.550 1.720 3.230 ;
        RECT  0.430 0.860 0.570 1.450 ;
        RECT  0.430 3.030 0.490 4.010 ;
        RECT  0.320 0.860 0.430 4.010 ;
        RECT  0.250 1.050 0.320 4.010 ;
        RECT  0.190 1.050 0.250 3.990 ;
        RECT  0.170 1.050 0.190 1.450 ;
    END
END SDFFTRX4

MACRO SDFFTRX2
    CLASS CORE ;
    FOREIGN SDFFTRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFTRXL ;
    SIZE 17.820 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.780 2.240 2.790 2.650 ;
        RECT  2.790 2.000 3.190 2.650 ;
        RECT  3.190 2.240 3.200 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.390 1.820 1.870 2.260 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.730 1.990 4.070 2.230 ;
        RECT  4.070 1.990 4.160 2.630 ;
        RECT  4.160 1.990 4.310 2.650 ;
        RECT  4.310 2.390 4.420 2.650 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.030 3.140 17.370 4.120 ;
        RECT  17.360 1.830 17.370 2.090 ;
        RECT  17.210 1.010 17.370 1.410 ;
        RECT  17.370 1.010 17.430 4.120 ;
        RECT  17.430 1.010 17.610 3.520 ;
        RECT  17.610 1.390 17.620 2.090 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.540 2.760 15.770 3.160 ;
        RECT  15.690 0.860 15.770 1.260 ;
        RECT  15.770 0.860 16.010 3.160 ;
        RECT  16.010 0.860 16.090 1.530 ;
        RECT  16.090 1.270 16.300 1.530 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.920 1.280 4.930 1.540 ;
        RECT  4.930 1.250 5.730 1.540 ;
        RECT  5.730 1.270 5.740 1.540 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.210 0.780 2.610 ;
        RECT  0.780 2.210 0.860 3.200 ;
        RECT  0.860 2.210 1.020 3.210 ;
        RECT  1.020 2.950 1.120 3.210 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.610 5.440 ;
        RECT  0.610 4.480 1.010 5.440 ;
        RECT  1.010 4.640 3.380 5.440 ;
        RECT  3.380 4.310 3.390 5.440 ;
        RECT  3.390 4.190 3.790 5.440 ;
        RECT  3.790 4.310 3.800 5.440 ;
        RECT  3.800 4.640 7.320 5.440 ;
        RECT  7.320 4.480 7.720 5.440 ;
        RECT  7.720 4.640 8.600 5.440 ;
        RECT  8.600 4.480 9.000 5.440 ;
        RECT  9.000 4.640 9.940 5.440 ;
        RECT  9.940 4.480 10.340 5.440 ;
        RECT  10.340 4.640 12.480 5.440 ;
        RECT  12.480 4.480 12.880 5.440 ;
        RECT  12.880 4.640 16.210 5.440 ;
        RECT  16.210 4.280 16.220 5.440 ;
        RECT  16.220 4.080 16.620 5.440 ;
        RECT  16.620 4.280 16.630 5.440 ;
        RECT  16.630 4.640 17.820 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.000 0.400 ;
        RECT  1.000 -0.400 1.010 1.350 ;
        RECT  1.010 -0.400 1.410 1.550 ;
        RECT  1.410 -0.400 1.420 1.350 ;
        RECT  1.420 -0.400 3.090 0.400 ;
        RECT  3.090 -0.400 3.490 0.560 ;
        RECT  3.490 -0.400 7.220 0.400 ;
        RECT  7.220 -0.400 7.230 0.730 ;
        RECT  7.230 -0.400 7.630 0.850 ;
        RECT  7.630 -0.400 7.640 0.730 ;
        RECT  7.640 -0.400 9.450 0.400 ;
        RECT  9.450 -0.400 9.460 0.840 ;
        RECT  9.460 -0.400 9.860 1.040 ;
        RECT  9.860 -0.400 9.870 0.840 ;
        RECT  9.870 -0.400 12.040 0.400 ;
        RECT  12.040 -0.400 12.050 0.980 ;
        RECT  12.050 -0.400 12.450 1.100 ;
        RECT  12.450 -0.400 12.460 0.980 ;
        RECT  12.460 -0.400 14.120 0.400 ;
        RECT  14.120 -0.400 14.130 1.100 ;
        RECT  14.130 -0.400 14.530 1.300 ;
        RECT  14.530 -0.400 14.540 1.100 ;
        RECT  14.540 -0.400 16.440 0.400 ;
        RECT  16.440 -0.400 16.450 0.690 ;
        RECT  16.450 -0.400 16.850 0.890 ;
        RECT  16.850 -0.400 16.860 0.690 ;
        RECT  16.860 -0.400 17.820 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.760 2.000 17.000 2.400 ;
        RECT  16.540 2.160 16.760 2.400 ;
        RECT  16.300 2.160 16.540 3.780 ;
        RECT  15.270 3.540 16.300 3.780 ;
        RECT  15.250 1.010 15.350 1.410 ;
        RECT  15.250 3.540 15.270 4.070 ;
        RECT  15.010 1.010 15.250 4.070 ;
        RECT  14.950 1.010 15.010 1.820 ;
        RECT  14.870 3.670 15.010 4.070 ;
        RECT  14.230 1.580 14.950 1.820 ;
        RECT  14.490 2.350 14.730 3.170 ;
        RECT  13.520 2.930 14.490 3.170 ;
        RECT  13.910 1.580 14.230 2.030 ;
        RECT  13.830 1.630 13.910 2.030 ;
        RECT  13.330 1.380 13.520 3.170 ;
        RECT  13.280 1.380 13.330 3.250 ;
        RECT  13.190 1.380 13.280 1.620 ;
        RECT  13.250 2.850 13.280 3.250 ;
        RECT  12.930 2.850 13.250 3.340 ;
        RECT  12.790 1.060 13.190 1.620 ;
        RECT  12.760 1.900 13.000 2.570 ;
        RECT  11.530 3.100 12.930 3.340 ;
        RECT  11.150 1.380 12.790 1.620 ;
        RECT  10.440 1.900 12.760 2.140 ;
        RECT  10.960 2.430 11.630 2.670 ;
        RECT  11.290 3.100 11.530 3.500 ;
        RECT  10.750 1.060 11.150 1.620 ;
        RECT  10.720 2.430 10.960 3.560 ;
        RECT  10.330 3.320 10.720 3.560 ;
        RECT  10.200 1.320 10.440 2.870 ;
        RECT  10.090 3.320 10.330 4.000 ;
        RECT  9.040 1.320 10.200 1.560 ;
        RECT  9.810 2.630 10.200 2.870 ;
        RECT  9.480 3.760 10.090 4.000 ;
        RECT  8.510 1.950 9.920 2.350 ;
        RECT  9.570 2.630 9.810 3.480 ;
        RECT  9.410 3.080 9.570 3.480 ;
        RECT  9.240 3.760 9.480 4.180 ;
        RECT  7.030 3.940 9.240 4.180 ;
        RECT  8.800 0.680 9.040 1.560 ;
        RECT  8.580 0.680 8.800 1.140 ;
        RECT  7.920 0.680 8.580 0.920 ;
        RECT  8.270 1.600 8.510 3.500 ;
        RECT  8.110 1.600 8.270 1.840 ;
        RECT  7.680 3.260 8.270 3.500 ;
        RECT  6.910 2.170 7.990 2.410 ;
        RECT  7.440 2.810 7.680 3.500 ;
        RECT  6.790 3.940 7.030 4.360 ;
        RECT  6.670 0.830 6.910 2.980 ;
        RECT  6.730 4.120 6.790 4.360 ;
        RECT  6.330 4.120 6.730 4.370 ;
        RECT  6.110 0.830 6.670 1.070 ;
        RECT  6.510 2.740 6.670 2.980 ;
        RECT  6.270 2.740 6.510 3.780 ;
        RECT  5.990 4.120 6.330 4.360 ;
        RECT  5.990 1.830 6.290 2.070 ;
        RECT  5.750 1.830 5.990 4.360 ;
        RECT  4.550 4.120 5.750 4.360 ;
        RECT  4.010 0.670 5.630 0.910 ;
        RECT  5.470 2.980 5.480 3.680 ;
        RECT  5.300 2.980 5.470 3.800 ;
        RECT  5.290 2.460 5.300 3.800 ;
        RECT  5.070 2.340 5.290 3.800 ;
        RECT  5.060 2.340 5.070 3.680 ;
        RECT  4.890 2.340 5.060 3.400 ;
        RECT  4.880 2.460 4.890 3.400 ;
        RECT  2.330 3.150 4.880 3.390 ;
        RECT  4.310 3.670 4.550 4.360 ;
        RECT  4.290 1.190 4.530 1.620 ;
        RECT  0.490 3.670 4.310 3.910 ;
        RECT  2.440 1.380 4.290 1.620 ;
        RECT  3.770 0.670 4.010 1.100 ;
        RECT  2.150 0.860 3.770 1.100 ;
        RECT  2.140 1.380 2.440 2.770 ;
        RECT  1.910 0.670 2.150 1.100 ;
        RECT  2.050 2.530 2.140 2.770 ;
        RECT  1.810 2.530 2.050 3.350 ;
        RECT  1.750 0.670 1.910 0.910 ;
        RECT  1.590 3.110 1.810 3.350 ;
        RECT  0.400 1.220 0.570 1.620 ;
        RECT  0.400 3.160 0.490 3.910 ;
        RECT  0.250 1.220 0.400 3.910 ;
        RECT  0.160 1.220 0.250 3.480 ;
    END
END SDFFTRX2

MACRO SDFFTRX1
    CLASS CORE ;
    FOREIGN SDFFTRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFTRXL ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.170 2.380 3.760 2.680 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.020 2.170 2.260 2.570 ;
        RECT  2.260 2.330 2.330 2.570 ;
        RECT  2.330 2.330 2.570 3.180 ;
        RECT  2.570 2.940 2.840 3.180 ;
        RECT  2.840 2.940 2.860 3.210 ;
        RECT  2.860 2.940 3.080 3.250 ;
        RECT  3.080 2.950 3.100 3.250 ;
        RECT  3.100 3.010 4.310 3.250 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.110 2.030 4.350 2.530 ;
        RECT  4.350 2.030 4.730 2.270 ;
        RECT  4.730 1.830 5.070 2.270 ;
        RECT  5.070 1.830 5.080 2.090 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.160 1.170 15.380 1.860 ;
        RECT  15.000 3.060 15.390 3.460 ;
        RECT  15.380 1.170 15.390 2.090 ;
        RECT  15.390 1.170 15.400 3.460 ;
        RECT  15.400 1.170 15.630 3.300 ;
        RECT  15.630 1.170 15.640 2.090 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.310 3.520 13.400 4.060 ;
        RECT  13.400 3.510 13.660 4.110 ;
        RECT  13.660 3.520 13.800 4.110 ;
        RECT  13.450 0.670 13.850 1.100 ;
        RECT  13.800 3.520 13.970 3.780 ;
        RECT  13.970 3.520 14.410 3.760 ;
        RECT  14.410 3.500 14.480 3.760 ;
        RECT  13.850 0.860 14.480 1.100 ;
        RECT  14.480 0.860 14.720 3.760 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.990 1.250 5.480 1.490 ;
        RECT  5.480 1.250 5.730 1.530 ;
        RECT  5.730 1.270 5.740 1.530 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.710 2.050 1.200 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.740 5.440 ;
        RECT  0.740 4.480 1.140 5.440 ;
        RECT  1.140 4.640 7.750 5.440 ;
        RECT  7.750 4.480 7.830 5.440 ;
        RECT  7.830 4.460 8.630 5.440 ;
        RECT  8.630 4.480 8.710 5.440 ;
        RECT  8.710 4.640 10.120 5.440 ;
        RECT  10.120 3.890 10.130 5.440 ;
        RECT  10.130 3.690 10.530 5.440 ;
        RECT  10.530 3.890 10.540 5.440 ;
        RECT  10.540 4.640 12.590 5.440 ;
        RECT  12.590 4.170 12.600 5.440 ;
        RECT  12.600 3.970 13.000 5.440 ;
        RECT  13.000 4.170 13.010 5.440 ;
        RECT  13.010 4.640 14.130 5.440 ;
        RECT  14.130 4.480 14.530 5.440 ;
        RECT  14.530 4.640 15.840 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.320 0.400 ;
        RECT  0.320 -0.400 0.720 0.560 ;
        RECT  0.720 -0.400 2.980 0.400 ;
        RECT  2.980 -0.400 3.380 0.560 ;
        RECT  3.380 -0.400 7.520 0.400 ;
        RECT  7.520 -0.400 7.530 0.950 ;
        RECT  7.530 -0.400 7.930 1.150 ;
        RECT  7.930 -0.400 7.940 0.950 ;
        RECT  7.940 -0.400 9.960 0.400 ;
        RECT  9.960 -0.400 9.970 1.130 ;
        RECT  9.970 -0.400 10.370 1.330 ;
        RECT  10.370 -0.400 10.380 1.130 ;
        RECT  10.380 -0.400 12.630 0.400 ;
        RECT  12.630 -0.400 13.030 0.560 ;
        RECT  13.030 -0.400 14.200 0.400 ;
        RECT  14.200 -0.400 14.600 0.560 ;
        RECT  14.600 -0.400 15.840 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  13.960 1.540 14.200 3.160 ;
        RECT  13.910 1.540 13.960 1.780 ;
        RECT  13.560 2.760 13.960 3.160 ;
        RECT  13.510 1.380 13.910 1.780 ;
        RECT  12.610 1.540 13.510 1.780 ;
        RECT  13.280 2.060 13.440 2.460 ;
        RECT  13.040 2.060 13.280 2.780 ;
        RECT  12.160 2.540 13.040 2.780 ;
        RECT  12.370 1.540 12.610 2.260 ;
        RECT  12.210 1.860 12.370 2.260 ;
        RECT  11.920 2.540 12.160 3.890 ;
        RECT  11.810 1.090 11.920 3.890 ;
        RECT  11.680 1.090 11.810 3.970 ;
        RECT  11.190 1.090 11.680 1.330 ;
        RECT  11.410 3.570 11.680 3.970 ;
        RECT  11.050 1.850 11.350 2.250 ;
        RECT  11.040 1.610 11.050 2.250 ;
        RECT  10.800 1.610 11.040 3.060 ;
        RECT  9.650 1.610 10.800 1.850 ;
        RECT  10.090 2.820 10.800 3.060 ;
        RECT  9.120 2.140 10.520 2.540 ;
        RECT  9.690 2.820 10.090 3.220 ;
        RECT  9.450 3.860 9.850 4.260 ;
        RECT  9.410 0.710 9.650 1.850 ;
        RECT  7.190 3.940 9.450 4.180 ;
        RECT  8.700 0.710 9.410 0.950 ;
        RECT  8.880 1.370 9.120 3.140 ;
        RECT  8.690 1.370 8.880 1.770 ;
        RECT  7.570 2.900 8.880 3.140 ;
        RECT  8.290 0.670 8.700 0.950 ;
        RECT  8.360 2.170 8.600 2.570 ;
        RECT  8.120 1.610 8.360 2.570 ;
        RECT  6.860 1.610 8.120 1.850 ;
        RECT  7.330 2.130 7.570 3.140 ;
        RECT  6.950 3.940 7.190 4.360 ;
        RECT  6.860 2.660 6.980 3.060 ;
        RECT  6.790 4.110 6.950 4.360 ;
        RECT  6.620 0.830 6.860 3.060 ;
        RECT  6.280 4.110 6.790 4.350 ;
        RECT  6.170 0.830 6.620 1.070 ;
        RECT  6.580 2.660 6.620 3.060 ;
        RECT  6.280 1.360 6.340 2.080 ;
        RECT  6.100 1.360 6.280 4.350 ;
        RECT  6.040 1.840 6.100 4.350 ;
        RECT  1.680 4.110 6.040 4.350 ;
        RECT  5.600 3.590 5.750 3.830 ;
        RECT  3.900 0.670 5.690 0.910 ;
        RECT  5.360 2.440 5.600 3.830 ;
        RECT  2.170 3.590 5.360 3.830 ;
        RECT  4.420 1.270 4.660 1.510 ;
        RECT  4.180 1.270 4.420 1.620 ;
        RECT  2.980 1.380 4.180 1.620 ;
        RECT  3.660 0.670 3.900 1.100 ;
        RECT  2.040 0.860 3.660 1.100 ;
        RECT  2.740 1.380 2.980 2.030 ;
        RECT  1.730 1.380 2.740 1.790 ;
        RECT  1.720 2.850 2.050 3.090 ;
        RECT  1.640 0.720 2.040 1.100 ;
        RECT  1.720 1.550 1.730 1.790 ;
        RECT  1.480 1.550 1.720 3.090 ;
        RECT  1.440 3.940 1.680 4.350 ;
        RECT  0.490 3.940 1.440 4.180 ;
        RECT  0.430 1.280 0.570 1.680 ;
        RECT  0.490 2.940 0.570 3.340 ;
        RECT  0.430 2.940 0.490 4.180 ;
        RECT  0.250 1.280 0.430 4.180 ;
        RECT  0.190 1.280 0.250 3.340 ;
        RECT  0.170 1.280 0.190 1.680 ;
        RECT  0.170 2.940 0.190 3.340 ;
    END
END SDFFTRX1

MACRO SDFFSRHQXL
    CLASS CORE ;
    FOREIGN SDFFSRHQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.460 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.720 4.130 9.490 4.370 ;
        RECT  9.490 3.570 9.730 4.370 ;
        RECT  9.730 3.570 10.530 3.810 ;
        RECT  10.530 3.570 10.770 4.370 ;
        RECT  10.770 4.130 13.290 4.370 ;
        RECT  13.290 3.660 13.530 4.370 ;
        RECT  13.530 3.660 13.650 3.900 ;
        RECT  13.650 3.520 13.750 3.900 ;
        RECT  13.750 3.500 13.930 3.900 ;
        RECT  13.930 2.390 14.170 3.900 ;
        RECT  14.170 2.390 14.370 2.700 ;
        RECT  14.370 2.460 14.450 2.700 ;
        RECT  14.170 3.660 17.790 3.900 ;
        RECT  17.590 2.340 17.790 2.580 ;
        RECT  17.790 2.340 18.030 3.900 ;
        RECT  18.030 2.640 18.270 2.960 ;
        RECT  18.270 2.640 18.370 2.940 ;
        RECT  18.370 2.700 18.950 2.940 ;
        RECT  18.950 2.620 19.350 3.020 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.250 2.390 3.650 2.790 ;
        RECT  3.650 2.390 3.750 2.710 ;
        RECT  3.750 2.390 3.760 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.740 1.280 4.820 2.300 ;
        RECT  4.820 1.270 4.980 2.300 ;
        RECT  4.980 1.270 5.080 1.530 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  16.210 2.390 16.700 2.630 ;
        RECT  16.700 2.390 16.960 2.650 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.660 3.420 19.060 3.820 ;
        RECT  19.060 3.420 19.250 3.780 ;
        RECT  19.250 3.420 19.350 3.760 ;
        RECT  19.350 3.420 19.720 3.660 ;
        RECT  18.820 1.260 19.720 1.540 ;
        RECT  19.720 1.260 19.960 3.660 ;
        RECT  19.960 1.260 19.970 1.540 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.950 1.690 3.210 ;
        RECT  1.690 2.170 1.780 3.210 ;
        RECT  1.780 2.170 1.930 3.200 ;
        RECT  1.930 2.170 2.210 2.570 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.740 2.230 0.770 2.650 ;
        RECT  0.770 2.220 1.210 2.660 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.880 5.440 ;
        RECT  0.880 4.480 1.280 5.440 ;
        RECT  1.280 4.640 2.690 5.440 ;
        RECT  2.690 4.280 2.700 5.440 ;
        RECT  2.700 4.160 3.100 5.440 ;
        RECT  3.100 4.280 3.110 5.440 ;
        RECT  3.110 4.640 7.040 5.440 ;
        RECT  7.040 4.480 7.440 5.440 ;
        RECT  7.440 4.640 10.010 5.440 ;
        RECT  10.010 4.090 10.250 5.440 ;
        RECT  10.250 4.640 13.800 5.440 ;
        RECT  13.800 4.300 13.810 5.440 ;
        RECT  13.810 4.180 14.210 5.440 ;
        RECT  14.210 4.300 14.220 5.440 ;
        RECT  14.220 4.640 15.700 5.440 ;
        RECT  15.700 4.480 16.100 5.440 ;
        RECT  16.100 4.640 17.380 5.440 ;
        RECT  17.380 4.480 17.780 5.440 ;
        RECT  17.780 4.640 19.480 5.440 ;
        RECT  19.480 4.480 19.880 5.440 ;
        RECT  19.880 4.640 20.460 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.440 0.400 ;
        RECT  0.440 -0.400 1.200 0.560 ;
        RECT  1.200 -0.400 3.010 0.400 ;
        RECT  3.010 -0.400 3.020 0.730 ;
        RECT  3.020 -0.400 3.420 0.850 ;
        RECT  3.420 -0.400 3.430 0.730 ;
        RECT  3.430 -0.400 6.910 0.400 ;
        RECT  6.910 -0.400 6.920 0.730 ;
        RECT  6.920 -0.400 7.320 0.930 ;
        RECT  7.320 -0.400 7.330 0.730 ;
        RECT  7.330 -0.400 10.600 0.400 ;
        RECT  10.600 -0.400 10.610 0.850 ;
        RECT  10.610 -0.400 11.010 0.970 ;
        RECT  11.010 -0.400 11.020 0.850 ;
        RECT  11.020 -0.400 13.540 0.400 ;
        RECT  13.540 -0.400 13.940 0.560 ;
        RECT  13.940 -0.400 17.300 0.400 ;
        RECT  17.300 -0.400 17.310 1.300 ;
        RECT  17.310 -0.400 17.710 1.500 ;
        RECT  17.710 -0.400 17.720 1.300 ;
        RECT  17.720 -0.400 20.460 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  18.470 0.750 20.050 0.990 ;
        RECT  19.030 1.820 19.430 2.300 ;
        RECT  16.830 1.820 19.030 2.060 ;
        RECT  18.230 0.750 18.470 1.540 ;
        RECT  18.070 1.140 18.230 1.540 ;
        RECT  16.860 3.080 17.510 3.320 ;
        RECT  16.540 2.960 16.860 3.320 ;
        RECT  16.430 1.320 16.830 2.060 ;
        RECT  15.100 0.670 16.690 0.910 ;
        RECT  15.920 2.960 16.540 3.200 ;
        RECT  15.920 1.820 16.430 2.060 ;
        RECT  15.680 1.820 15.920 3.200 ;
        RECT  15.380 2.250 15.680 2.650 ;
        RECT  14.980 1.460 15.400 1.700 ;
        RECT  14.780 0.670 15.100 1.130 ;
        RECT  14.740 1.460 14.980 3.380 ;
        RECT  13.070 0.890 14.780 1.130 ;
        RECT  13.650 1.460 14.740 1.700 ;
        RECT  14.500 2.980 14.740 3.380 ;
        RECT  13.410 1.460 13.650 2.760 ;
        RECT  12.830 0.890 13.070 3.270 ;
        RECT  12.610 3.540 13.010 3.850 ;
        RECT  12.310 0.890 12.830 1.130 ;
        RECT  12.260 3.030 12.830 3.270 ;
        RECT  11.260 3.540 12.610 3.810 ;
        RECT  12.310 1.410 12.550 2.690 ;
        RECT  11.810 1.410 12.310 1.650 ;
        RECT  11.900 2.450 12.310 2.690 ;
        RECT  11.290 1.930 12.030 2.170 ;
        RECT  11.580 2.450 11.900 3.250 ;
        RECT  11.570 1.250 11.810 1.650 ;
        RECT  11.500 2.890 11.580 3.250 ;
        RECT  11.260 1.250 11.290 2.170 ;
        RECT  11.050 1.250 11.260 3.810 ;
        RECT  9.970 1.250 11.050 1.490 ;
        RECT  11.020 1.930 11.050 3.810 ;
        RECT  11.010 2.930 11.020 3.810 ;
        RECT  9.860 2.930 11.010 3.170 ;
        RECT  10.530 1.770 10.770 2.570 ;
        RECT  8.690 1.770 10.530 2.010 ;
        RECT  9.730 0.670 9.970 1.490 ;
        RECT  9.210 2.290 9.760 2.530 ;
        RECT  9.560 0.670 9.730 0.910 ;
        RECT  8.970 2.290 9.210 3.850 ;
        RECT  6.710 3.610 8.970 3.850 ;
        RECT  8.450 1.270 8.690 3.330 ;
        RECT  8.410 1.270 8.450 1.670 ;
        RECT  7.090 3.090 8.450 3.330 ;
        RECT  7.930 2.000 8.170 2.410 ;
        RECT  6.300 2.000 7.930 2.240 ;
        RECT  6.850 2.520 7.090 3.330 ;
        RECT  6.690 2.520 6.850 2.760 ;
        RECT  6.470 3.610 6.710 4.350 ;
        RECT  5.500 4.110 6.470 4.350 ;
        RECT  6.060 0.910 6.300 2.740 ;
        RECT  5.670 0.910 6.060 1.310 ;
        RECT  6.020 2.500 6.060 2.740 ;
        RECT  5.780 2.500 6.020 3.820 ;
        RECT  5.500 1.820 5.780 2.060 ;
        RECT  5.260 1.820 5.500 4.350 ;
        RECT  3.620 4.110 5.260 4.350 ;
        RECT  3.940 0.670 5.190 0.910 ;
        RECT  4.140 3.590 4.980 3.830 ;
        RECT  4.480 2.600 4.720 3.170 ;
        RECT  4.460 2.600 4.480 2.840 ;
        RECT  4.220 1.330 4.460 2.840 ;
        RECT  2.930 1.650 4.220 1.890 ;
        RECT  3.900 3.120 4.140 3.830 ;
        RECT  3.700 0.670 3.940 1.370 ;
        RECT  2.210 3.120 3.900 3.360 ;
        RECT  2.140 1.130 3.700 1.370 ;
        RECT  3.380 3.640 3.620 4.350 ;
        RECT  0.490 3.640 3.380 3.880 ;
        RECT  2.530 1.650 2.930 2.720 ;
        RECT  1.410 1.650 2.530 1.890 ;
        RECT  1.170 1.530 1.410 1.930 ;
        RECT  0.450 1.390 0.850 1.790 ;
        RECT  0.450 2.930 0.490 3.880 ;
        RECT  0.250 1.390 0.450 3.880 ;
        RECT  0.210 1.390 0.250 3.230 ;
    END
END SDFFSRHQXL

MACRO SDFFSRHQX4
    CLASS CORE ;
    FOREIGN SDFFSRHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSRHQXL ;
    SIZE 28.380 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.880 4.130 10.180 4.370 ;
        RECT  10.180 3.660 10.420 4.370 ;
        RECT  10.420 3.660 10.450 4.200 ;
        RECT  10.450 3.660 13.310 3.900 ;
        RECT  13.310 3.660 13.550 4.370 ;
        RECT  13.550 4.130 16.880 4.370 ;
        RECT  16.880 3.660 17.120 4.370 ;
        RECT  17.120 3.660 17.340 3.900 ;
        RECT  17.340 2.380 17.710 3.900 ;
        RECT  17.710 2.380 17.740 2.780 ;
        RECT  17.710 3.660 20.770 3.900 ;
        RECT  20.770 3.020 21.010 3.900 ;
        RECT  21.010 3.020 25.430 3.260 ;
        RECT  25.430 2.340 25.670 3.260 ;
        RECT  25.670 2.340 26.240 2.580 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.430 2.250 3.840 2.790 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.890 1.260 4.900 1.540 ;
        RECT  4.900 1.260 5.140 2.270 ;
        RECT  5.140 1.260 5.740 1.540 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  19.820 2.320 19.920 2.720 ;
        RECT  19.920 2.310 20.520 2.730 ;
        RECT  20.520 2.320 20.800 2.720 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.710 3.540 22.110 3.940 ;
        RECT  22.150 1.310 22.550 1.710 ;
        RECT  22.550 1.390 23.860 1.630 ;
        RECT  22.110 3.540 24.150 3.780 ;
        RECT  23.860 1.310 24.260 1.710 ;
        RECT  24.150 3.540 24.750 3.940 ;
        RECT  24.260 1.390 25.390 1.630 ;
        RECT  25.390 1.310 25.550 1.710 ;
        RECT  25.550 1.310 25.790 2.060 ;
        RECT  25.790 1.820 26.070 2.060 ;
        RECT  24.750 3.540 26.130 3.780 ;
        RECT  26.130 3.000 26.510 3.980 ;
        RECT  26.070 1.820 26.510 2.100 ;
        RECT  26.510 1.820 26.530 3.980 ;
        RECT  26.530 1.820 26.930 3.410 ;
        RECT  26.930 1.820 26.950 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.380 1.990 2.660 ;
        RECT  1.990 2.170 2.390 2.660 ;
        RECT  2.390 2.380 2.400 2.660 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.690 2.340 0.720 2.740 ;
        RECT  0.720 2.340 1.070 3.220 ;
        RECT  1.070 2.340 1.110 3.210 ;
        RECT  1.110 2.950 1.120 3.210 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 4.480 1.390 5.440 ;
        RECT  1.390 4.640 2.850 5.440 ;
        RECT  2.850 4.280 2.860 5.440 ;
        RECT  2.860 4.160 3.260 5.440 ;
        RECT  3.260 4.280 3.270 5.440 ;
        RECT  3.270 4.640 7.200 5.440 ;
        RECT  7.200 4.480 7.600 5.440 ;
        RECT  7.600 4.640 10.690 5.440 ;
        RECT  10.690 4.310 10.700 5.440 ;
        RECT  10.700 4.190 11.100 5.440 ;
        RECT  11.100 4.310 11.110 5.440 ;
        RECT  11.110 4.640 12.390 5.440 ;
        RECT  12.390 4.300 12.400 5.440 ;
        RECT  12.400 4.180 12.800 5.440 ;
        RECT  12.800 4.300 12.810 5.440 ;
        RECT  12.810 4.640 17.390 5.440 ;
        RECT  17.390 4.300 17.400 5.440 ;
        RECT  17.400 4.180 17.800 5.440 ;
        RECT  17.800 4.300 17.810 5.440 ;
        RECT  17.810 4.640 19.240 5.440 ;
        RECT  19.240 4.480 19.640 5.440 ;
        RECT  19.640 4.640 20.910 5.440 ;
        RECT  20.910 4.480 21.310 5.440 ;
        RECT  21.310 4.640 22.920 5.440 ;
        RECT  22.920 4.320 22.930 5.440 ;
        RECT  22.930 4.120 23.330 5.440 ;
        RECT  23.330 4.320 23.340 5.440 ;
        RECT  23.340 4.640 25.360 5.440 ;
        RECT  25.360 4.320 25.370 5.440 ;
        RECT  25.370 4.120 25.770 5.440 ;
        RECT  25.770 4.320 25.780 5.440 ;
        RECT  25.780 4.640 26.880 5.440 ;
        RECT  26.880 4.160 26.890 5.440 ;
        RECT  26.890 3.960 27.290 5.440 ;
        RECT  27.290 4.160 27.300 5.440 ;
        RECT  27.300 4.640 28.380 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.920 0.400 ;
        RECT  0.920 -0.400 0.930 1.060 ;
        RECT  0.930 -0.400 1.330 1.260 ;
        RECT  1.330 -0.400 1.340 1.060 ;
        RECT  1.340 -0.400 3.110 0.400 ;
        RECT  3.110 -0.400 3.120 0.730 ;
        RECT  3.120 -0.400 3.520 0.850 ;
        RECT  3.520 -0.400 3.530 0.730 ;
        RECT  3.530 -0.400 7.010 0.400 ;
        RECT  7.010 -0.400 7.250 0.930 ;
        RECT  7.250 -0.400 10.880 0.400 ;
        RECT  10.880 -0.400 10.890 0.980 ;
        RECT  10.890 -0.400 11.290 1.100 ;
        RECT  11.290 -0.400 11.300 0.980 ;
        RECT  11.300 -0.400 12.460 0.400 ;
        RECT  12.460 -0.400 12.470 1.110 ;
        RECT  12.470 -0.400 12.870 1.230 ;
        RECT  12.870 -0.400 12.880 1.110 ;
        RECT  12.880 -0.400 16.650 0.400 ;
        RECT  16.650 -0.400 17.050 0.560 ;
        RECT  17.050 -0.400 20.510 0.400 ;
        RECT  20.510 -0.400 20.520 1.120 ;
        RECT  20.520 -0.400 20.920 1.320 ;
        RECT  20.920 -0.400 20.930 1.120 ;
        RECT  20.930 -0.400 27.040 0.400 ;
        RECT  27.040 -0.400 27.050 0.800 ;
        RECT  27.050 -0.400 27.450 1.000 ;
        RECT  27.450 -0.400 27.460 0.800 ;
        RECT  27.460 -0.400 28.380 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  27.730 1.280 28.130 1.680 ;
        RECT  26.310 1.280 27.730 1.520 ;
        RECT  26.070 0.750 26.310 1.520 ;
        RECT  25.110 0.750 26.070 0.990 ;
        RECT  24.710 0.670 25.110 1.070 ;
        RECT  24.670 1.960 25.070 2.360 ;
        RECT  23.280 0.750 24.710 0.990 ;
        RECT  24.650 2.040 24.670 2.360 ;
        RECT  23.310 2.040 24.650 2.280 ;
        RECT  23.300 2.040 23.310 2.540 ;
        RECT  22.900 2.040 23.300 2.730 ;
        RECT  22.880 0.670 23.280 1.070 ;
        RECT  22.890 2.040 22.900 2.540 ;
        RECT  21.640 2.040 22.890 2.280 ;
        RECT  21.400 1.320 21.640 2.280 ;
        RECT  21.240 1.320 21.400 2.010 ;
        RECT  20.200 1.770 21.240 2.010 ;
        RECT  19.250 3.080 20.490 3.320 ;
        RECT  19.800 1.320 20.200 2.010 ;
        RECT  18.310 0.730 19.850 0.970 ;
        RECT  19.250 1.770 19.800 2.010 ;
        RECT  19.010 1.770 19.250 3.320 ;
        RECT  18.280 1.460 18.620 1.700 ;
        RECT  17.990 0.730 18.310 1.120 ;
        RECT  18.040 1.460 18.280 3.380 ;
        RECT  16.780 1.460 18.040 1.700 ;
        RECT  17.990 2.980 18.040 3.380 ;
        RECT  17.910 0.860 17.990 1.120 ;
        RECT  15.820 0.860 17.910 1.100 ;
        RECT  16.540 1.460 16.780 2.240 ;
        RECT  16.340 3.560 16.600 3.800 ;
        RECT  16.100 3.560 16.340 3.850 ;
        RECT  15.750 2.880 16.270 3.280 ;
        RECT  14.110 3.610 16.100 3.850 ;
        RECT  15.750 0.860 15.820 1.570 ;
        RECT  15.660 0.860 15.750 3.330 ;
        RECT  15.510 0.670 15.660 3.330 ;
        RECT  15.420 0.670 15.510 1.570 ;
        RECT  14.390 3.090 15.510 3.330 ;
        RECT  14.380 0.670 15.420 0.910 ;
        RECT  14.940 1.250 15.100 1.490 ;
        RECT  14.700 1.250 14.940 1.750 ;
        RECT  14.350 1.510 14.700 1.750 ;
        RECT  14.140 0.670 14.380 1.230 ;
        RECT  14.110 1.510 14.350 2.800 ;
        RECT  13.980 0.990 14.140 1.230 ;
        RECT  13.630 1.510 14.110 1.750 ;
        RECT  13.760 2.560 14.110 2.800 ;
        RECT  13.870 3.140 14.110 3.850 ;
        RECT  11.300 3.140 13.870 3.380 ;
        RECT  11.300 2.030 13.830 2.270 ;
        RECT  13.440 2.560 13.760 2.860 ;
        RECT  13.230 1.170 13.630 1.750 ;
        RECT  11.580 2.620 13.440 2.860 ;
        RECT  12.110 1.510 13.230 1.750 ;
        RECT  11.710 1.170 12.110 1.750 ;
        RECT  11.060 1.380 11.300 3.380 ;
        RECT  10.420 1.380 11.060 1.620 ;
        RECT  10.200 3.000 11.060 3.240 ;
        RECT  10.520 1.900 10.760 2.570 ;
        RECT  9.360 1.900 10.520 2.140 ;
        RECT  10.000 0.660 10.420 1.630 ;
        RECT  9.880 2.420 10.120 2.660 ;
        RECT  9.710 0.670 10.000 0.910 ;
        RECT  9.640 2.420 9.880 3.850 ;
        RECT  9.430 1.220 9.670 1.620 ;
        RECT  6.710 3.610 9.640 3.850 ;
        RECT  9.190 0.750 9.430 1.620 ;
        RECT  9.120 1.900 9.360 3.230 ;
        RECT  8.150 0.750 9.190 0.990 ;
        RECT  8.910 1.900 9.120 2.140 ;
        RECT  7.250 2.990 9.120 3.230 ;
        RECT  8.650 1.270 8.910 2.140 ;
        RECT  8.140 2.420 8.690 2.660 ;
        RECT  8.510 1.270 8.650 1.670 ;
        RECT  7.910 0.750 8.150 1.630 ;
        RECT  7.900 2.000 8.140 2.660 ;
        RECT  7.750 1.230 7.910 1.630 ;
        RECT  6.660 2.000 7.900 2.240 ;
        RECT  7.010 2.520 7.250 3.230 ;
        RECT  6.790 2.520 7.010 2.760 ;
        RECT  6.470 3.610 6.710 4.350 ;
        RECT  6.460 0.750 6.660 2.240 ;
        RECT  5.660 4.110 6.470 4.350 ;
        RECT  6.220 0.750 6.460 2.740 ;
        RECT  5.750 0.750 6.220 0.990 ;
        RECT  6.180 2.500 6.220 2.740 ;
        RECT  5.940 2.500 6.180 3.550 ;
        RECT  5.660 1.820 5.940 2.060 ;
        RECT  5.420 1.820 5.660 4.350 ;
        RECT  3.780 4.110 5.420 4.350 ;
        RECT  4.040 0.750 5.390 0.990 ;
        RECT  4.300 3.590 5.140 3.830 ;
        RECT  4.660 2.550 4.900 3.170 ;
        RECT  4.560 2.550 4.660 2.790 ;
        RECT  4.320 1.330 4.560 2.790 ;
        RECT  3.110 1.650 4.320 1.890 ;
        RECT  4.060 3.070 4.300 3.830 ;
        RECT  2.370 3.070 4.060 3.310 ;
        RECT  3.800 0.750 4.040 1.370 ;
        RECT  2.240 1.130 3.800 1.370 ;
        RECT  3.540 3.640 3.780 4.350 ;
        RECT  0.570 3.640 3.540 3.880 ;
        RECT  2.710 1.650 3.110 2.720 ;
        RECT  1.680 1.650 2.710 1.890 ;
        RECT  1.280 1.650 1.680 1.940 ;
        RECT  0.410 1.120 0.570 1.520 ;
        RECT  0.410 3.490 0.570 3.890 ;
        RECT  0.170 1.120 0.410 3.890 ;
    END
END SDFFSRHQX4

MACRO SDFFSRHQX2
    CLASS CORE ;
    FOREIGN SDFFSRHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSRHQXL ;
    SIZE 24.420 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.720 4.130 9.490 4.370 ;
        RECT  9.490 3.660 9.730 4.370 ;
        RECT  9.730 3.660 12.750 3.900 ;
        RECT  12.750 3.660 12.920 4.080 ;
        RECT  12.920 3.660 13.160 4.370 ;
        RECT  13.160 4.130 16.400 4.370 ;
        RECT  16.400 3.660 16.640 4.370 ;
        RECT  16.700 2.950 16.800 3.210 ;
        RECT  16.640 3.660 16.810 3.900 ;
        RECT  16.800 2.540 16.810 3.210 ;
        RECT  16.810 2.540 16.900 3.900 ;
        RECT  16.900 2.380 17.050 3.900 ;
        RECT  17.050 2.380 17.300 2.780 ;
        RECT  17.050 3.660 18.210 3.900 ;
        RECT  18.210 3.610 18.450 3.900 ;
        RECT  18.450 3.610 20.650 3.850 ;
        RECT  20.650 3.020 20.890 3.850 ;
        RECT  20.890 3.020 22.230 3.260 ;
        RECT  22.230 2.940 22.380 3.260 ;
        RECT  22.380 2.770 22.770 3.260 ;
        RECT  22.770 2.770 23.150 3.010 ;
        RECT  23.150 2.040 23.160 3.010 ;
        RECT  23.160 1.960 23.390 3.010 ;
        RECT  23.390 1.960 23.560 2.360 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.260 2.390 3.660 2.790 ;
        RECT  3.660 2.390 3.750 2.710 ;
        RECT  3.750 2.390 3.760 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.740 1.280 4.820 2.300 ;
        RECT  4.820 1.270 4.980 2.300 ;
        RECT  4.980 1.270 5.080 1.530 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  19.250 2.310 19.850 2.730 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.740 3.540 22.140 3.940 ;
        RECT  22.140 3.540 22.770 3.780 ;
        RECT  22.770 3.500 23.210 3.780 ;
        RECT  23.210 3.500 23.840 3.790 ;
        RECT  21.930 1.390 23.840 1.630 ;
        RECT  23.840 1.390 24.080 3.980 ;
        RECT  24.080 3.000 24.240 3.980 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.160 2.230 2.650 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.740 2.070 0.770 2.470 ;
        RECT  0.770 1.820 1.110 2.470 ;
        RECT  1.110 1.820 1.120 2.120 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.880 5.440 ;
        RECT  0.880 4.480 1.280 5.440 ;
        RECT  1.280 4.640 2.690 5.440 ;
        RECT  2.690 4.280 2.700 5.440 ;
        RECT  2.700 4.160 3.100 5.440 ;
        RECT  3.100 4.280 3.110 5.440 ;
        RECT  3.110 4.640 7.040 5.440 ;
        RECT  7.040 4.480 7.440 5.440 ;
        RECT  7.440 4.640 10.000 5.440 ;
        RECT  10.000 4.300 10.010 5.440 ;
        RECT  10.010 4.180 10.410 5.440 ;
        RECT  10.410 4.300 10.420 5.440 ;
        RECT  10.420 4.640 12.010 5.440 ;
        RECT  12.010 4.300 12.020 5.440 ;
        RECT  12.020 4.180 12.420 5.440 ;
        RECT  12.420 4.300 12.430 5.440 ;
        RECT  12.430 4.640 16.910 5.440 ;
        RECT  16.910 4.300 16.920 5.440 ;
        RECT  16.920 4.180 17.320 5.440 ;
        RECT  17.320 4.300 17.330 5.440 ;
        RECT  17.330 4.640 18.850 5.440 ;
        RECT  18.850 4.480 19.250 5.440 ;
        RECT  19.250 4.640 20.440 5.440 ;
        RECT  20.440 4.480 20.840 5.440 ;
        RECT  20.840 4.640 23.070 5.440 ;
        RECT  23.070 4.370 23.080 5.440 ;
        RECT  23.080 4.250 23.480 5.440 ;
        RECT  23.480 4.370 23.490 5.440 ;
        RECT  23.490 4.640 24.420 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.280 0.400 ;
        RECT  0.280 -0.400 0.680 0.560 ;
        RECT  0.680 -0.400 3.010 0.400 ;
        RECT  3.010 -0.400 3.020 0.730 ;
        RECT  3.020 -0.400 3.420 0.850 ;
        RECT  3.420 -0.400 3.430 0.730 ;
        RECT  3.430 -0.400 6.780 0.400 ;
        RECT  6.780 -0.400 6.790 0.730 ;
        RECT  6.790 -0.400 7.190 0.850 ;
        RECT  7.190 -0.400 7.200 0.730 ;
        RECT  7.200 -0.400 10.600 0.400 ;
        RECT  10.600 -0.400 10.610 0.730 ;
        RECT  10.610 -0.400 11.010 0.850 ;
        RECT  11.010 -0.400 11.020 0.730 ;
        RECT  11.020 -0.400 12.100 0.400 ;
        RECT  12.100 -0.400 12.110 1.110 ;
        RECT  12.110 -0.400 12.510 1.230 ;
        RECT  12.510 -0.400 12.520 1.110 ;
        RECT  12.520 -0.400 16.440 0.400 ;
        RECT  16.440 -0.400 16.840 0.560 ;
        RECT  16.840 -0.400 20.200 0.400 ;
        RECT  20.200 -0.400 20.210 1.120 ;
        RECT  20.210 -0.400 20.610 1.320 ;
        RECT  20.610 -0.400 20.620 1.120 ;
        RECT  20.620 -0.400 23.840 0.400 ;
        RECT  23.840 -0.400 23.850 0.670 ;
        RECT  23.850 -0.400 24.250 0.870 ;
        RECT  24.250 -0.400 24.260 0.670 ;
        RECT  24.260 -0.400 24.420 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  21.540 0.790 23.240 1.030 ;
        RECT  22.410 1.960 22.810 2.360 ;
        RECT  20.750 2.040 22.410 2.280 ;
        RECT  21.140 0.670 21.540 1.030 ;
        RECT  20.510 1.770 20.750 2.280 ;
        RECT  19.840 1.770 20.510 2.010 ;
        RECT  18.860 3.080 20.100 3.320 ;
        RECT  19.440 1.320 19.840 2.010 ;
        RECT  17.960 0.670 19.500 0.910 ;
        RECT  18.860 1.770 19.440 2.010 ;
        RECT  18.620 1.770 18.860 3.320 ;
        RECT  17.840 1.460 18.270 1.700 ;
        RECT  17.640 0.670 17.960 1.120 ;
        RECT  17.840 2.990 17.920 3.300 ;
        RECT  17.600 1.460 17.840 3.300 ;
        RECT  17.560 0.860 17.640 1.120 ;
        RECT  16.510 1.460 17.600 1.700 ;
        RECT  17.520 2.990 17.600 3.300 ;
        RECT  15.550 0.860 17.560 1.100 ;
        RECT  16.270 1.460 16.510 2.240 ;
        RECT  13.750 3.610 16.120 3.850 ;
        RECT  15.390 2.930 15.770 3.330 ;
        RECT  15.390 0.860 15.550 1.580 ;
        RECT  15.150 0.670 15.390 3.330 ;
        RECT  14.050 0.670 15.150 0.910 ;
        RECT  14.030 3.090 15.150 3.330 ;
        RECT  14.640 1.250 14.800 1.490 ;
        RECT  14.400 1.250 14.640 1.750 ;
        RECT  13.990 1.510 14.400 1.750 ;
        RECT  13.810 0.670 14.050 1.230 ;
        RECT  13.750 1.510 13.990 2.800 ;
        RECT  13.640 0.990 13.810 1.230 ;
        RECT  13.270 1.510 13.750 1.750 ;
        RECT  13.220 2.560 13.750 2.800 ;
        RECT  13.510 3.140 13.750 3.850 ;
        RECT  10.940 3.140 13.510 3.380 ;
        RECT  10.940 2.030 13.470 2.270 ;
        RECT  12.870 1.170 13.270 1.750 ;
        RECT  12.900 2.560 13.220 2.860 ;
        RECT  11.220 2.620 12.900 2.860 ;
        RECT  11.750 1.510 12.870 1.750 ;
        RECT  11.350 1.170 11.750 1.750 ;
        RECT  10.700 1.250 10.940 3.380 ;
        RECT  9.970 1.250 10.700 1.490 ;
        RECT  9.860 2.930 10.700 3.170 ;
        RECT  10.160 1.770 10.400 2.570 ;
        RECT  8.690 1.770 10.160 2.010 ;
        RECT  9.730 0.670 9.970 1.490 ;
        RECT  9.210 2.290 9.760 2.530 ;
        RECT  9.560 0.670 9.730 0.910 ;
        RECT  8.970 2.290 9.210 3.850 ;
        RECT  6.710 3.610 8.970 3.850 ;
        RECT  8.450 1.270 8.690 3.330 ;
        RECT  8.410 1.270 8.450 1.670 ;
        RECT  7.090 3.090 8.450 3.330 ;
        RECT  7.930 2.000 8.170 2.410 ;
        RECT  6.300 2.000 7.930 2.240 ;
        RECT  6.850 2.520 7.090 3.330 ;
        RECT  6.690 2.520 6.850 2.760 ;
        RECT  6.470 3.610 6.710 4.350 ;
        RECT  5.500 4.110 6.470 4.350 ;
        RECT  6.060 0.990 6.300 2.740 ;
        RECT  5.670 0.990 6.060 1.230 ;
        RECT  6.020 2.500 6.060 2.740 ;
        RECT  5.780 2.500 6.020 3.830 ;
        RECT  5.500 1.820 5.780 2.060 ;
        RECT  5.260 1.820 5.500 4.350 ;
        RECT  3.620 4.110 5.260 4.350 ;
        RECT  3.940 0.670 5.190 0.910 ;
        RECT  4.140 3.590 4.980 3.830 ;
        RECT  4.490 2.600 4.730 3.170 ;
        RECT  4.460 2.600 4.490 2.840 ;
        RECT  4.220 1.330 4.460 2.840 ;
        RECT  2.940 1.650 4.220 1.890 ;
        RECT  3.900 3.120 4.140 3.830 ;
        RECT  3.700 0.670 3.940 1.370 ;
        RECT  2.210 3.120 3.900 3.360 ;
        RECT  2.140 1.130 3.700 1.370 ;
        RECT  3.380 3.640 3.620 4.350 ;
        RECT  0.570 3.640 3.380 3.880 ;
        RECT  2.540 1.650 2.940 2.720 ;
        RECT  1.860 1.650 2.540 1.890 ;
        RECT  1.620 0.640 1.860 1.890 ;
        RECT  1.460 0.640 1.620 0.880 ;
        RECT  0.450 3.070 0.570 3.880 ;
        RECT  0.450 1.390 0.490 1.790 ;
        RECT  0.330 1.390 0.450 3.880 ;
        RECT  0.210 1.390 0.330 3.470 ;
        RECT  0.170 3.070 0.210 3.470 ;
    END
END SDFFSRHQX2

MACRO SDFFSRHQX1
    CLASS CORE ;
    FOREIGN SDFFSRHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSRHQXL ;
    SIZE 20.460 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.720 4.130 9.490 4.370 ;
        RECT  9.490 3.570 9.730 4.370 ;
        RECT  9.730 3.570 10.530 3.810 ;
        RECT  10.530 3.570 10.770 4.370 ;
        RECT  10.770 4.130 13.290 4.370 ;
        RECT  13.290 3.660 13.530 4.370 ;
        RECT  13.530 3.660 13.650 3.900 ;
        RECT  13.650 3.520 13.750 3.900 ;
        RECT  13.750 3.500 13.930 3.900 ;
        RECT  13.930 2.390 14.170 3.900 ;
        RECT  14.170 2.390 14.370 2.700 ;
        RECT  14.370 2.460 14.450 2.700 ;
        RECT  14.170 3.660 17.790 3.900 ;
        RECT  17.590 2.340 17.790 2.580 ;
        RECT  17.790 2.340 18.030 3.900 ;
        RECT  18.030 2.640 18.270 2.960 ;
        RECT  18.270 2.640 18.370 2.940 ;
        RECT  18.370 2.700 18.950 2.940 ;
        RECT  18.950 2.620 19.350 3.020 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.250 2.390 3.650 2.790 ;
        RECT  3.650 2.390 3.750 2.710 ;
        RECT  3.750 2.390 3.760 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.740 1.280 4.820 2.300 ;
        RECT  4.820 1.270 4.980 2.300 ;
        RECT  4.980 1.270 5.080 1.530 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  16.210 2.400 16.700 2.640 ;
        RECT  16.700 2.390 16.960 2.650 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.660 3.630 19.060 4.030 ;
        RECT  18.710 1.280 19.340 1.520 ;
        RECT  19.060 3.630 19.590 3.870 ;
        RECT  19.340 1.270 19.600 1.530 ;
        RECT  19.590 3.520 19.630 3.870 ;
        RECT  19.600 1.290 19.630 1.530 ;
        RECT  19.630 1.290 19.870 3.870 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.390 1.630 2.650 ;
        RECT  1.630 2.320 2.030 2.720 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.740 2.070 0.770 2.470 ;
        RECT  0.770 1.830 1.110 2.470 ;
        RECT  1.110 1.830 1.130 2.120 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.880 5.440 ;
        RECT  0.880 4.480 1.280 5.440 ;
        RECT  1.280 4.640 2.690 5.440 ;
        RECT  2.690 4.280 2.700 5.440 ;
        RECT  2.700 4.160 3.100 5.440 ;
        RECT  3.100 4.280 3.110 5.440 ;
        RECT  3.110 4.640 7.040 5.440 ;
        RECT  7.040 4.480 7.440 5.440 ;
        RECT  7.440 4.640 10.010 5.440 ;
        RECT  10.010 4.090 10.250 5.440 ;
        RECT  10.250 4.640 13.800 5.440 ;
        RECT  13.800 4.300 13.810 5.440 ;
        RECT  13.810 4.180 14.210 5.440 ;
        RECT  14.210 4.300 14.220 5.440 ;
        RECT  14.220 4.640 15.750 5.440 ;
        RECT  15.750 4.480 16.150 5.440 ;
        RECT  16.150 4.640 17.380 5.440 ;
        RECT  17.380 4.480 17.780 5.440 ;
        RECT  17.780 4.640 19.480 5.440 ;
        RECT  19.480 4.480 19.880 5.440 ;
        RECT  19.880 4.640 20.460 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.310 0.400 ;
        RECT  0.310 -0.400 0.710 0.560 ;
        RECT  0.710 -0.400 3.010 0.400 ;
        RECT  3.010 -0.400 3.020 0.730 ;
        RECT  3.020 -0.400 3.420 0.850 ;
        RECT  3.420 -0.400 3.430 0.730 ;
        RECT  3.430 -0.400 6.910 0.400 ;
        RECT  6.910 -0.400 6.920 0.730 ;
        RECT  6.920 -0.400 7.320 0.850 ;
        RECT  7.320 -0.400 7.330 0.730 ;
        RECT  7.330 -0.400 10.600 0.400 ;
        RECT  10.600 -0.400 10.610 0.730 ;
        RECT  10.610 -0.400 11.010 0.850 ;
        RECT  11.010 -0.400 11.020 0.730 ;
        RECT  11.020 -0.400 13.540 0.400 ;
        RECT  13.540 -0.400 13.940 0.560 ;
        RECT  13.940 -0.400 17.180 0.400 ;
        RECT  17.180 -0.400 17.190 1.420 ;
        RECT  17.190 -0.400 17.590 1.540 ;
        RECT  17.590 -0.400 17.600 1.420 ;
        RECT  17.600 -0.400 20.460 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  18.350 0.750 19.930 0.990 ;
        RECT  19.270 1.980 19.350 2.220 ;
        RECT  18.950 1.820 19.270 2.220 ;
        RECT  16.750 1.820 18.950 2.060 ;
        RECT  18.110 0.750 18.350 1.460 ;
        RECT  17.950 1.060 18.110 1.460 ;
        RECT  15.920 3.080 17.510 3.320 ;
        RECT  16.510 1.320 16.750 2.060 ;
        RECT  15.100 0.670 16.630 0.910 ;
        RECT  15.920 1.820 16.510 2.060 ;
        RECT  15.680 1.820 15.920 3.320 ;
        RECT  15.520 2.250 15.680 2.650 ;
        RECT  14.980 1.460 15.400 1.700 ;
        RECT  14.780 0.670 15.100 1.120 ;
        RECT  14.740 1.460 14.980 3.380 ;
        RECT  14.700 0.860 14.780 1.120 ;
        RECT  13.650 1.460 14.740 1.700 ;
        RECT  14.500 2.980 14.740 3.380 ;
        RECT  13.070 0.860 14.700 1.100 ;
        RECT  13.410 1.460 13.650 2.760 ;
        RECT  12.830 0.860 13.070 3.270 ;
        RECT  12.610 3.570 13.010 3.850 ;
        RECT  12.310 0.890 12.830 1.130 ;
        RECT  12.260 3.030 12.830 3.270 ;
        RECT  11.340 3.570 12.610 3.810 ;
        RECT  12.310 1.410 12.550 2.690 ;
        RECT  11.810 1.410 12.310 1.650 ;
        RECT  11.820 2.450 12.310 2.690 ;
        RECT  11.340 1.930 12.030 2.170 ;
        RECT  11.580 2.450 11.820 3.330 ;
        RECT  11.570 1.250 11.810 1.650 ;
        RECT  11.290 1.930 11.340 3.810 ;
        RECT  11.100 1.130 11.290 3.810 ;
        RECT  11.050 1.130 11.100 2.170 ;
        RECT  9.860 2.930 11.100 3.170 ;
        RECT  10.130 1.130 11.050 1.370 ;
        RECT  10.530 1.770 10.770 2.570 ;
        RECT  8.690 1.770 10.530 2.010 ;
        RECT  9.970 1.130 10.130 1.490 ;
        RECT  9.730 0.670 9.970 1.490 ;
        RECT  9.210 2.290 9.760 2.530 ;
        RECT  9.560 0.670 9.730 0.910 ;
        RECT  8.970 2.290 9.210 3.850 ;
        RECT  6.710 3.610 8.970 3.850 ;
        RECT  8.450 1.270 8.690 3.330 ;
        RECT  8.410 1.270 8.450 1.670 ;
        RECT  7.090 3.090 8.450 3.330 ;
        RECT  7.930 2.000 8.170 2.410 ;
        RECT  6.300 2.000 7.930 2.240 ;
        RECT  6.850 2.520 7.090 3.330 ;
        RECT  6.690 2.520 6.850 2.760 ;
        RECT  6.470 3.610 6.710 4.350 ;
        RECT  5.500 4.110 6.470 4.350 ;
        RECT  6.060 0.990 6.300 2.740 ;
        RECT  5.670 0.990 6.060 1.230 ;
        RECT  6.020 2.500 6.060 2.740 ;
        RECT  5.780 2.500 6.020 3.830 ;
        RECT  5.500 1.820 5.780 2.060 ;
        RECT  5.260 1.820 5.500 4.350 ;
        RECT  3.620 4.110 5.260 4.350 ;
        RECT  3.940 0.670 5.190 0.910 ;
        RECT  4.140 3.590 4.980 3.830 ;
        RECT  4.480 2.600 4.720 3.170 ;
        RECT  4.460 2.600 4.480 2.840 ;
        RECT  4.220 1.330 4.460 2.840 ;
        RECT  2.910 1.650 4.220 1.890 ;
        RECT  3.900 3.120 4.140 3.830 ;
        RECT  3.700 0.670 3.940 1.370 ;
        RECT  2.210 3.120 3.900 3.360 ;
        RECT  2.140 1.130 3.700 1.370 ;
        RECT  3.380 3.640 3.620 4.350 ;
        RECT  0.490 3.640 3.380 3.880 ;
        RECT  2.510 1.650 2.910 2.720 ;
        RECT  2.500 1.650 2.510 2.640 ;
        RECT  1.860 1.650 2.500 1.890 ;
        RECT  1.620 0.680 1.860 1.890 ;
        RECT  1.460 0.680 1.620 0.920 ;
        RECT  0.450 1.390 0.490 1.790 ;
        RECT  0.450 2.840 0.490 3.880 ;
        RECT  0.250 1.390 0.450 3.880 ;
        RECT  0.210 1.390 0.250 3.230 ;
    END
END SDFFSRHQX1

MACRO SDFFSRXL
    CLASS CORE ;
    FOREIGN SDFFSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.150 3.940 7.550 4.370 ;
        RECT  7.550 3.940 8.530 4.180 ;
        RECT  8.530 3.940 8.770 4.360 ;
        RECT  8.770 4.080 8.790 4.360 ;
        RECT  8.790 4.120 10.420 4.360 ;
        RECT  10.420 4.120 10.770 4.370 ;
        RECT  10.770 4.130 14.060 4.370 ;
        RECT  14.060 4.070 14.070 4.370 ;
        RECT  14.070 4.030 14.310 4.370 ;
        RECT  14.310 4.030 14.320 4.330 ;
        RECT  14.320 4.030 14.730 4.270 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.950 2.850 3.210 ;
        RECT  2.850 2.190 3.090 3.210 ;
        RECT  3.090 2.950 3.100 3.210 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.950 0.210 3.210 ;
        RECT  0.210 2.560 0.460 3.210 ;
        RECT  0.460 2.560 0.530 3.200 ;
        RECT  0.530 2.560 0.610 2.960 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.120 1.270 8.270 1.530 ;
        RECT  8.270 1.270 8.380 1.950 ;
        RECT  8.380 1.280 8.510 1.950 ;
        RECT  8.510 1.710 8.710 1.950 ;
        RECT  8.710 1.710 8.950 2.110 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.700 2.950 16.900 3.210 ;
        RECT  16.800 1.390 16.900 1.790 ;
        RECT  16.900 1.390 17.140 3.240 ;
        RECT  17.140 1.390 17.200 1.790 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.020 2.950 18.030 3.210 ;
        RECT  18.030 2.840 18.690 3.240 ;
        RECT  18.570 1.350 18.690 1.750 ;
        RECT  18.690 2.640 18.730 3.240 ;
        RECT  18.690 1.350 18.730 1.840 ;
        RECT  18.730 1.350 18.970 3.240 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.720 2.190 2.120 2.630 ;
        RECT  2.120 2.390 2.180 2.630 ;
        RECT  2.180 2.390 2.440 2.650 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  10.620 2.360 11.220 2.710 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.370 5.440 ;
        RECT  0.370 4.480 0.770 5.440 ;
        RECT  0.770 4.640 3.310 5.440 ;
        RECT  3.310 4.480 3.710 5.440 ;
        RECT  3.710 4.640 6.250 5.440 ;
        RECT  6.250 4.480 6.650 5.440 ;
        RECT  6.650 4.640 7.850 5.440 ;
        RECT  7.850 4.480 8.250 5.440 ;
        RECT  11.170 3.520 11.570 3.850 ;
        RECT  11.570 3.610 13.460 3.850 ;
        RECT  13.460 3.360 13.700 3.850 ;
        RECT  8.250 4.640 15.060 5.440 ;
        RECT  13.700 3.360 15.060 3.600 ;
        RECT  15.060 3.360 15.300 5.440 ;
        RECT  15.300 4.640 15.900 5.440 ;
        RECT  15.900 3.700 15.910 5.440 ;
        RECT  15.910 3.580 16.310 5.440 ;
        RECT  16.310 3.700 16.320 5.440 ;
        RECT  16.320 4.640 17.630 5.440 ;
        RECT  17.630 4.480 18.030 5.440 ;
        RECT  18.030 4.640 19.140 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.470 0.400 ;
        RECT  0.470 -0.400 0.480 1.490 ;
        RECT  0.480 -0.400 0.790 1.710 ;
        RECT  0.790 1.470 0.880 1.710 ;
        RECT  0.790 -0.400 3.280 0.400 ;
        RECT  3.280 -0.400 3.680 0.560 ;
        RECT  3.680 -0.400 5.870 0.400 ;
        RECT  5.870 -0.400 5.880 0.730 ;
        RECT  5.880 -0.400 6.280 0.850 ;
        RECT  6.280 -0.400 6.290 0.730 ;
        RECT  6.290 -0.400 9.300 0.400 ;
        RECT  9.300 -0.400 9.310 0.730 ;
        RECT  9.310 -0.400 9.710 0.850 ;
        RECT  9.710 -0.400 9.720 0.730 ;
        RECT  9.720 -0.400 11.200 0.400 ;
        RECT  11.200 -0.400 11.210 1.450 ;
        RECT  11.210 -0.400 11.610 1.570 ;
        RECT  11.610 -0.400 11.620 1.450 ;
        RECT  11.620 -0.400 13.830 0.400 ;
        RECT  13.830 -0.400 13.840 1.290 ;
        RECT  13.840 -0.400 14.240 1.490 ;
        RECT  14.240 -0.400 14.250 1.290 ;
        RECT  14.250 -0.400 17.680 0.400 ;
        RECT  17.680 -0.400 18.080 0.560 ;
        RECT  18.080 -0.400 19.140 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  18.270 2.030 18.450 2.430 ;
        RECT  18.030 0.860 18.270 2.430 ;
        RECT  17.200 0.860 18.030 1.100 ;
        RECT  17.660 2.190 18.030 2.430 ;
        RECT  17.420 2.190 17.660 3.910 ;
        RECT  17.160 3.670 17.420 3.910 ;
        RECT  16.800 0.730 17.200 1.100 ;
        RECT  16.760 3.670 17.160 4.070 ;
        RECT  15.860 2.190 16.620 2.590 ;
        RECT  15.620 1.260 15.860 3.080 ;
        RECT  15.380 1.260 15.620 1.500 ;
        RECT  13.890 2.840 15.620 3.080 ;
        RECT  13.180 2.210 15.330 2.450 ;
        RECT  13.490 2.790 13.890 3.080 ;
        RECT  12.170 0.680 13.220 0.920 ;
        RECT  12.940 1.330 13.180 3.330 ;
        RECT  12.500 1.330 12.940 1.570 ;
        RECT  12.450 3.090 12.940 3.330 ;
        RECT  12.170 2.520 12.550 2.760 ;
        RECT  11.930 0.680 12.170 3.220 ;
        RECT  10.730 1.850 11.930 2.090 ;
        RECT  10.730 2.980 11.930 3.220 ;
        RECT  10.490 1.650 10.730 2.090 ;
        RECT  10.490 2.980 10.730 3.840 ;
        RECT  10.420 0.780 10.580 1.020 ;
        RECT  10.320 1.650 10.490 1.890 ;
        RECT  9.290 3.600 10.490 3.840 ;
        RECT  10.180 0.780 10.420 1.370 ;
        RECT  9.030 1.130 10.180 1.370 ;
        RECT  9.740 2.430 9.970 3.320 ;
        RECT  9.630 2.420 9.740 3.320 ;
        RECT  9.570 1.650 9.630 3.320 ;
        RECT  9.390 1.650 9.570 3.140 ;
        RECT  9.220 1.650 9.390 1.890 ;
        RECT  8.510 2.900 9.390 3.140 ;
        RECT  9.050 3.420 9.290 3.840 ;
        RECT  5.730 3.420 9.050 3.660 ;
        RECT  8.790 0.750 9.030 1.370 ;
        RECT  7.760 0.750 8.790 0.990 ;
        RECT  8.270 2.430 8.510 3.140 ;
        RECT  7.760 1.810 7.990 3.140 ;
        RECT  7.750 0.750 7.760 3.140 ;
        RECT  7.520 0.750 7.750 2.050 ;
        RECT  6.230 2.900 7.750 3.140 ;
        RECT  7.240 2.330 7.470 2.570 ;
        RECT  7.000 1.130 7.240 2.570 ;
        RECT  5.710 1.130 7.000 1.370 ;
        RECT  5.990 2.740 6.230 3.140 ;
        RECT  5.490 3.420 5.730 4.370 ;
        RECT  5.470 1.130 5.710 3.120 ;
        RECT  5.330 4.130 5.490 4.370 ;
        RECT  5.160 1.130 5.470 1.370 ;
        RECT  5.190 2.880 5.470 3.120 ;
        RECT  4.960 1.880 5.190 2.280 ;
        RECT  4.950 2.880 5.190 3.290 ;
        RECT  4.830 0.720 5.160 1.370 ;
        RECT  4.400 1.880 4.960 2.290 ;
        RECT  4.760 0.720 4.830 0.960 ;
        RECT  4.400 3.250 4.620 3.650 ;
        RECT  4.020 0.720 4.420 1.100 ;
        RECT  4.160 1.470 4.400 3.650 ;
        RECT  4.130 3.940 4.370 4.370 ;
        RECT  3.840 1.470 4.160 1.710 ;
        RECT  3.730 3.230 4.160 3.650 ;
        RECT  3.260 3.940 4.130 4.180 ;
        RECT  2.250 0.860 4.020 1.100 ;
        RECT  3.020 3.610 3.260 4.180 ;
        RECT  2.250 3.610 3.020 3.850 ;
        RECT  1.320 4.130 2.470 4.370 ;
        RECT  1.840 0.670 2.250 1.100 ;
        RECT  2.010 3.200 2.250 3.850 ;
        RECT  1.850 3.200 2.010 3.440 ;
        RECT  1.430 0.670 1.510 0.910 ;
        RECT  1.320 0.670 1.430 2.320 ;
        RECT  1.190 0.670 1.320 4.370 ;
        RECT  1.110 0.670 1.190 0.910 ;
        RECT  1.080 2.000 1.190 4.370 ;
    END
END SDFFSRXL

MACRO SDFFSRX4
    CLASS CORE ;
    FOREIGN SDFFSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSRXL ;
    SIZE 25.740 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.420 3.990 7.820 4.360 ;
        RECT  7.820 4.120 11.310 4.360 ;
        RECT  11.310 3.940 11.760 4.360 ;
        RECT  11.760 3.940 16.170 4.180 ;
        RECT  16.170 3.940 16.870 4.340 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.950 2.900 3.210 ;
        RECT  2.900 2.150 3.100 3.210 ;
        RECT  3.100 2.150 3.140 3.200 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.700 2.380 1.200 2.840 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.360 2.380 9.900 2.810 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  23.000 2.750 23.210 3.150 ;
        RECT  23.190 1.390 23.210 1.790 ;
        RECT  23.210 1.390 23.610 3.220 ;
        RECT  23.610 1.820 23.650 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  24.530 1.390 24.930 3.220 ;
        RECT  24.930 1.820 24.970 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.810 2.580 2.180 2.820 ;
        RECT  2.180 2.390 2.430 2.820 ;
        RECT  2.430 2.390 2.440 2.650 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.760 2.090 ;
        RECT  3.760 1.850 4.000 2.350 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.780 5.440 ;
        RECT  0.780 4.480 1.180 5.440 ;
        RECT  1.180 4.640 3.120 5.440 ;
        RECT  3.120 4.480 3.520 5.440 ;
        RECT  3.520 4.640 6.740 5.440 ;
        RECT  6.740 4.480 7.140 5.440 ;
        RECT  7.140 4.640 12.250 5.440 ;
        RECT  12.250 4.480 12.650 5.440 ;
        RECT  12.650 4.640 14.780 5.440 ;
        RECT  14.780 4.480 15.180 5.440 ;
        RECT  15.180 4.640 17.710 5.440 ;
        RECT  17.710 3.100 18.110 5.440 ;
        RECT  18.110 4.640 19.610 5.440 ;
        RECT  19.610 3.610 20.010 5.440 ;
        RECT  20.010 4.640 22.360 5.440 ;
        RECT  22.360 4.010 22.760 5.440 ;
        RECT  22.760 4.640 23.760 5.440 ;
        RECT  23.760 4.210 23.770 5.440 ;
        RECT  23.770 4.010 24.170 5.440 ;
        RECT  24.170 4.210 24.180 5.440 ;
        RECT  24.180 4.640 25.180 5.440 ;
        RECT  25.180 4.010 25.580 5.440 ;
        RECT  25.580 4.640 25.740 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.820 0.400 ;
        RECT  0.820 -0.400 0.830 0.730 ;
        RECT  0.830 -0.400 1.230 0.930 ;
        RECT  1.230 -0.400 1.240 0.730 ;
        RECT  1.240 -0.400 3.340 0.400 ;
        RECT  3.340 -0.400 3.740 0.560 ;
        RECT  3.740 -0.400 6.520 0.400 ;
        RECT  6.520 -0.400 6.530 0.730 ;
        RECT  6.530 -0.400 6.930 0.850 ;
        RECT  6.930 -0.400 6.940 0.730 ;
        RECT  6.940 -0.400 9.340 0.400 ;
        RECT  9.340 -0.400 9.350 0.800 ;
        RECT  9.350 -0.400 9.750 0.920 ;
        RECT  9.750 -0.400 9.760 0.800 ;
        RECT  9.760 -0.400 12.230 0.400 ;
        RECT  12.230 -0.400 12.470 1.400 ;
        RECT  12.470 -0.400 14.640 0.400 ;
        RECT  14.640 -0.400 14.650 0.820 ;
        RECT  14.650 -0.400 15.050 0.940 ;
        RECT  15.050 -0.400 15.060 0.820 ;
        RECT  15.060 -0.400 17.580 0.400 ;
        RECT  17.580 -0.400 17.590 0.880 ;
        RECT  17.590 -0.400 17.990 1.080 ;
        RECT  17.990 -0.400 18.000 0.880 ;
        RECT  18.000 -0.400 22.540 0.400 ;
        RECT  22.540 -0.400 22.550 0.910 ;
        RECT  22.550 -0.400 22.950 1.110 ;
        RECT  22.950 -0.400 22.960 0.910 ;
        RECT  22.960 -0.400 23.850 0.400 ;
        RECT  23.850 -0.400 23.860 0.910 ;
        RECT  23.860 -0.400 24.260 1.110 ;
        RECT  24.260 -0.400 24.270 0.910 ;
        RECT  24.270 -0.400 25.160 0.400 ;
        RECT  25.160 -0.400 25.170 0.910 ;
        RECT  25.170 -0.400 25.570 1.110 ;
        RECT  25.570 -0.400 25.580 0.910 ;
        RECT  25.580 -0.400 25.740 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  25.210 2.170 25.450 3.730 ;
        RECT  22.760 3.490 25.210 3.730 ;
        RECT  22.520 1.550 22.760 3.730 ;
        RECT  22.050 1.550 22.520 1.790 ;
        RECT  21.510 3.330 22.520 3.730 ;
        RECT  21.880 2.130 22.280 2.530 ;
        RECT  21.810 1.390 22.050 1.790 ;
        RECT  21.570 2.140 21.880 2.530 ;
        RECT  20.200 0.720 21.620 0.960 ;
        RECT  21.330 1.480 21.570 3.050 ;
        RECT  20.920 1.480 21.330 1.720 ;
        RECT  21.190 2.810 21.330 3.050 ;
        RECT  20.950 2.810 21.190 3.640 ;
        RECT  20.810 2.060 21.050 2.460 ;
        RECT  20.790 3.080 20.950 3.640 ;
        RECT  20.500 1.200 20.920 1.720 ;
        RECT  18.940 2.060 20.810 2.300 ;
        RECT  18.830 3.080 20.790 3.320 ;
        RECT  19.460 1.480 20.500 1.720 ;
        RECT  19.780 0.720 20.200 1.200 ;
        RECT  18.740 0.720 19.780 0.960 ;
        RECT  19.220 1.240 19.460 1.720 ;
        RECT  19.060 1.240 19.220 1.480 ;
        RECT  18.700 1.920 18.940 2.300 ;
        RECT  18.670 3.080 18.830 3.630 ;
        RECT  18.580 0.720 18.740 1.320 ;
        RECT  16.600 1.920 18.700 2.160 ;
        RECT  18.430 2.580 18.670 3.630 ;
        RECT  18.500 0.720 18.580 1.610 ;
        RECT  18.340 0.920 18.500 1.610 ;
        RECT  17.390 2.580 18.430 2.820 ;
        RECT  17.150 1.370 18.340 1.610 ;
        RECT  17.230 3.420 17.470 4.370 ;
        RECT  17.150 2.580 17.390 3.100 ;
        RECT  11.180 3.420 17.230 3.660 ;
        RECT  16.910 0.940 17.150 1.610 ;
        RECT  15.480 2.860 17.150 3.100 ;
        RECT  16.360 0.830 16.600 2.160 ;
        RECT  15.990 0.830 16.360 1.070 ;
        RECT  16.120 1.920 16.360 2.160 ;
        RECT  15.720 1.920 16.120 2.620 ;
        RECT  14.930 1.400 16.070 1.640 ;
        RECT  14.210 1.920 15.720 2.160 ;
        RECT  15.240 2.440 15.480 3.100 ;
        RECT  15.080 2.440 15.240 2.680 ;
        RECT  14.690 1.220 14.930 1.640 ;
        RECT  14.230 1.220 14.690 1.460 ;
        RECT  13.990 0.670 14.230 1.460 ;
        RECT  13.970 1.750 14.210 3.140 ;
        RECT  13.170 0.670 13.990 0.910 ;
        RECT  13.690 1.750 13.970 1.990 ;
        RECT  13.520 2.900 13.970 3.140 ;
        RECT  13.450 1.190 13.690 1.990 ;
        RECT  13.170 2.270 13.690 2.510 ;
        RECT  12.930 0.670 13.170 2.510 ;
        RECT  12.360 2.270 12.930 2.510 ;
        RECT  12.120 2.040 12.360 2.510 ;
        RECT  11.950 2.040 12.120 2.280 ;
        RECT  11.680 2.900 11.840 3.140 ;
        RECT  11.650 2.560 11.680 3.140 ;
        RECT  11.440 1.370 11.650 3.140 ;
        RECT  10.400 0.770 11.530 1.010 ;
        RECT  11.410 1.370 11.440 2.800 ;
        RECT  10.810 2.020 11.410 2.260 ;
        RECT  10.940 3.080 11.180 3.660 ;
        RECT  10.470 3.080 10.940 3.320 ;
        RECT  8.340 3.600 10.660 3.840 ;
        RECT  10.230 1.720 10.470 3.320 ;
        RECT  10.160 0.770 10.400 1.440 ;
        RECT  10.050 1.720 10.230 1.960 ;
        RECT  9.030 3.080 10.230 3.320 ;
        RECT  8.510 1.200 10.160 1.440 ;
        RECT  8.790 2.370 9.030 3.320 ;
        RECT  8.270 1.200 8.510 3.100 ;
        RECT  8.100 3.470 8.340 3.840 ;
        RECT  8.010 1.200 8.270 1.440 ;
        RECT  8.090 2.860 8.270 3.100 ;
        RECT  6.330 3.470 8.100 3.710 ;
        RECT  7.690 2.860 8.090 3.190 ;
        RECT  7.690 1.770 7.930 2.270 ;
        RECT  5.870 1.770 7.690 2.010 ;
        RECT  6.710 2.860 7.690 3.100 ;
        RECT  6.470 2.300 6.710 3.100 ;
        RECT  6.090 3.470 6.330 4.330 ;
        RECT  5.270 4.090 6.090 4.330 ;
        RECT  5.800 0.670 5.870 2.010 ;
        RECT  5.790 0.670 5.800 2.420 ;
        RECT  5.560 0.670 5.790 3.820 ;
        RECT  5.410 0.670 5.560 0.910 ;
        RECT  5.550 2.180 5.560 3.820 ;
        RECT  4.620 1.490 5.280 1.890 ;
        RECT  5.030 3.210 5.270 4.330 ;
        RECT  4.810 0.670 5.050 0.910 ;
        RECT  4.620 3.210 5.030 3.450 ;
        RECT  4.570 0.670 4.810 1.100 ;
        RECT  4.510 3.730 4.750 4.130 ;
        RECT  4.380 1.410 4.620 3.450 ;
        RECT  2.610 0.860 4.570 1.100 ;
        RECT  3.590 3.730 4.510 3.970 ;
        RECT  4.210 1.410 4.380 1.650 ;
        RECT  3.930 2.990 4.380 3.450 ;
        RECT  3.350 3.490 3.590 3.970 ;
        RECT  2.450 3.490 3.350 3.730 ;
        RECT  1.690 4.010 2.710 4.250 ;
        RECT  2.370 0.860 2.610 1.650 ;
        RECT  2.050 3.100 2.450 3.730 ;
        RECT  2.210 1.250 2.370 1.650 ;
        RECT  1.450 3.180 1.690 4.250 ;
        RECT  0.570 1.860 1.590 2.100 ;
        RECT  0.410 3.180 1.450 3.420 ;
        RECT  0.410 1.370 0.570 2.100 ;
        RECT  0.170 1.370 0.410 3.420 ;
    END
END SDFFSRX4

MACRO SDFFSRX2
    CLASS CORE ;
    FOREIGN SDFFSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSRXL ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.530 3.940 6.930 4.370 ;
        RECT  6.930 3.940 8.030 4.180 ;
        RECT  8.030 3.940 8.270 4.360 ;
        RECT  8.270 4.120 10.210 4.360 ;
        RECT  10.210 4.120 10.450 4.370 ;
        RECT  10.450 4.130 13.650 4.370 ;
        RECT  13.650 4.080 13.800 4.370 ;
        RECT  13.800 4.030 14.200 4.370 ;
        RECT  14.200 4.030 14.310 4.330 ;
        RECT  14.310 4.070 14.320 4.330 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.600 2.350 2.750 2.750 ;
        RECT  2.750 2.350 2.760 2.940 ;
        RECT  2.760 2.350 2.840 3.200 ;
        RECT  2.840 2.350 3.000 3.210 ;
        RECT  3.000 2.950 3.100 3.210 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.660 2.680 0.860 3.200 ;
        RECT  0.860 2.680 0.900 3.210 ;
        RECT  0.900 2.950 1.120 3.210 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.120 1.830 8.130 2.090 ;
        RECT  8.130 1.780 8.760 2.180 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.140 1.160 17.220 1.560 ;
        RECT  17.220 1.160 17.460 3.210 ;
        RECT  17.460 1.160 17.540 1.560 ;
        RECT  17.460 2.950 17.620 3.210 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.580 3.180 18.690 4.160 ;
        RECT  18.690 2.950 18.730 4.160 ;
        RECT  18.580 1.020 18.730 1.420 ;
        RECT  18.730 1.020 18.970 4.160 ;
        RECT  18.970 3.180 18.980 4.160 ;
        RECT  18.970 1.020 18.980 1.420 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.330 2.250 1.870 2.660 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  10.100 2.250 10.850 2.720 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 3.080 5.440 ;
        RECT  3.080 4.480 3.480 5.440 ;
        RECT  3.480 4.640 5.860 5.440 ;
        RECT  5.860 4.480 6.260 5.440 ;
        RECT  6.260 4.640 7.390 5.440 ;
        RECT  7.390 4.480 7.790 5.440 ;
        RECT  10.890 3.510 11.290 3.850 ;
        RECT  11.290 3.610 13.100 3.850 ;
        RECT  13.100 3.460 13.340 3.850 ;
        RECT  7.790 4.640 14.710 5.440 ;
        RECT  13.340 3.460 14.710 3.700 ;
        RECT  14.710 3.460 14.950 5.440 ;
        RECT  14.950 4.640 15.620 5.440 ;
        RECT  15.620 3.730 15.630 5.440 ;
        RECT  15.630 3.530 16.030 5.440 ;
        RECT  16.030 3.730 16.040 5.440 ;
        RECT  16.040 4.640 17.860 5.440 ;
        RECT  17.860 4.150 18.260 5.440 ;
        RECT  18.260 4.640 19.140 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.440 0.400 ;
        RECT  0.440 -0.400 0.840 0.950 ;
        RECT  0.840 -0.400 2.890 0.400 ;
        RECT  2.890 -0.400 3.290 0.560 ;
        RECT  3.290 -0.400 5.870 0.400 ;
        RECT  5.870 -0.400 5.880 0.730 ;
        RECT  5.880 -0.400 6.280 0.930 ;
        RECT  6.280 -0.400 6.290 0.730 ;
        RECT  6.290 -0.400 8.950 0.400 ;
        RECT  8.950 -0.400 9.350 0.850 ;
        RECT  9.350 -0.400 10.990 0.400 ;
        RECT  10.990 -0.400 11.390 1.410 ;
        RECT  11.390 -0.400 13.310 0.400 ;
        RECT  13.310 -0.400 13.710 0.560 ;
        RECT  13.710 -0.400 16.360 0.400 ;
        RECT  16.360 -0.400 16.760 0.560 ;
        RECT  16.760 -0.400 17.860 0.400 ;
        RECT  17.860 -0.400 18.260 1.710 ;
        RECT  18.260 -0.400 19.140 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  18.290 2.320 18.490 2.560 ;
        RECT  18.050 2.320 18.290 3.830 ;
        RECT  16.900 3.590 18.050 3.830 ;
        RECT  16.820 1.290 16.900 3.830 ;
        RECT  16.760 1.290 16.820 3.990 ;
        RECT  16.660 1.130 16.760 3.990 ;
        RECT  16.360 1.130 16.660 1.530 ;
        RECT  16.420 3.590 16.660 3.990 ;
        RECT  16.180 1.820 16.420 3.170 ;
        RECT  15.300 1.820 16.180 2.060 ;
        RECT  13.600 2.930 16.180 3.170 ;
        RECT  15.540 0.750 15.940 1.150 ;
        RECT  14.500 0.750 15.540 0.990 ;
        RECT  15.060 1.270 15.300 2.060 ;
        RECT  14.820 1.270 15.060 1.510 ;
        RECT  14.580 1.850 14.820 2.260 ;
        RECT  12.710 1.850 14.580 2.090 ;
        RECT  14.100 0.750 14.500 1.150 ;
        RECT  13.360 2.610 13.600 3.170 ;
        RECT  13.190 2.610 13.360 2.850 ;
        RECT  11.940 0.730 12.930 0.970 ;
        RECT  12.580 1.410 12.710 3.330 ;
        RECT  12.470 1.250 12.580 3.330 ;
        RECT  12.180 1.250 12.470 1.650 ;
        RECT  12.190 3.090 12.470 3.330 ;
        RECT  11.940 2.520 12.230 2.760 ;
        RECT  11.700 0.730 11.940 3.230 ;
        RECT  10.510 1.740 11.700 1.980 ;
        RECT  10.450 2.990 11.700 3.230 ;
        RECT  10.110 1.360 10.510 1.980 ;
        RECT  10.210 2.990 10.450 3.880 ;
        RECT  9.830 0.770 10.370 1.010 ;
        RECT  8.750 3.640 10.210 3.880 ;
        RECT  9.590 0.770 9.830 1.370 ;
        RECT  9.390 2.430 9.680 2.830 ;
        RECT  7.820 1.130 9.590 1.370 ;
        RECT  9.390 1.650 9.440 1.890 ;
        RECT  9.150 1.650 9.390 3.390 ;
        RECT  9.040 1.650 9.150 1.890 ;
        RECT  8.990 2.900 9.150 3.390 ;
        RECT  8.260 2.900 8.990 3.140 ;
        RECT  8.510 3.420 8.750 3.880 ;
        RECT  5.550 3.420 8.510 3.660 ;
        RECT  8.020 2.510 8.260 3.140 ;
        RECT  7.740 1.110 7.820 1.510 ;
        RECT  7.500 1.110 7.740 3.140 ;
        RECT  7.420 1.110 7.500 1.510 ;
        RECT  6.060 2.900 7.500 3.140 ;
        RECT  6.980 1.810 7.220 2.210 ;
        RECT  5.540 1.970 6.980 2.210 ;
        RECT  5.820 2.490 6.060 3.140 ;
        RECT  5.310 3.420 5.550 4.370 ;
        RECT  5.300 1.030 5.540 2.970 ;
        RECT  5.050 4.130 5.310 4.370 ;
        RECT  4.960 1.030 5.300 1.270 ;
        RECT  5.020 2.730 5.300 2.970 ;
        RECT  4.780 1.740 5.020 2.140 ;
        RECT  4.780 2.730 5.020 3.850 ;
        RECT  4.560 0.870 4.960 1.270 ;
        RECT  4.370 1.740 4.780 1.980 ;
        RECT  4.370 3.250 4.450 3.650 ;
        RECT  4.130 1.740 4.370 3.650 ;
        RECT  3.900 3.940 4.140 4.360 ;
        RECT  4.030 1.740 4.130 1.980 ;
        RECT  3.560 3.300 4.130 3.650 ;
        RECT  3.630 0.670 4.030 1.100 ;
        RECT  3.630 1.390 4.030 1.980 ;
        RECT  3.260 3.940 3.900 4.180 ;
        RECT  2.260 0.860 3.630 1.100 ;
        RECT  3.020 3.610 3.260 4.180 ;
        RECT  2.020 3.610 3.020 3.850 ;
        RECT  2.020 0.860 2.260 1.590 ;
        RECT  1.090 4.130 2.240 4.370 ;
        RECT  1.950 1.350 2.020 1.590 ;
        RECT  1.620 3.310 2.020 3.850 ;
        RECT  1.710 1.350 1.950 1.750 ;
        RECT  1.360 0.640 1.730 0.880 ;
        RECT  1.120 0.640 1.360 1.630 ;
        RECT  1.010 1.390 1.120 1.630 ;
        RECT  0.850 3.940 1.090 4.370 ;
        RECT  0.770 1.390 1.010 2.360 ;
        RECT  0.380 3.940 0.850 4.180 ;
        RECT  0.610 1.960 0.770 2.360 ;
        RECT  0.380 2.120 0.610 2.360 ;
        RECT  0.140 2.120 0.380 4.180 ;
    END
END SDFFSRX2

MACRO SDFFSRX1
    CLASS CORE ;
    FOREIGN SDFFSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSRXL ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.570 3.940 6.970 4.350 ;
        RECT  6.970 3.940 7.950 4.180 ;
        RECT  7.950 3.940 8.190 4.360 ;
        RECT  8.190 4.120 10.110 4.360 ;
        RECT  10.110 4.120 10.350 4.370 ;
        RECT  10.350 4.130 13.650 4.370 ;
        RECT  13.650 4.080 13.700 4.370 ;
        RECT  13.700 4.030 14.310 4.370 ;
        RECT  14.310 4.070 14.320 4.330 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.600 2.350 2.750 2.750 ;
        RECT  2.750 2.350 2.760 2.940 ;
        RECT  2.760 2.350 2.840 3.190 ;
        RECT  2.840 2.350 3.000 3.210 ;
        RECT  3.000 2.950 3.100 3.210 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.680 0.860 3.200 ;
        RECT  0.860 2.680 0.920 3.210 ;
        RECT  0.920 2.950 1.120 3.210 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.110 1.820 8.520 2.190 ;
        RECT  8.520 1.780 8.760 2.190 ;
        RECT  8.760 1.820 8.770 2.190 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.390 0.730 16.630 3.750 ;
        RECT  16.630 3.510 16.700 3.750 ;
        RECT  16.700 3.510 16.880 3.770 ;
        RECT  16.880 3.510 17.120 4.150 ;
        RECT  17.120 3.750 17.290 4.150 ;
        RECT  16.630 0.730 17.290 0.970 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.020 2.950 18.130 3.210 ;
        RECT  18.130 2.940 18.530 3.220 ;
        RECT  18.530 2.940 18.660 3.430 ;
        RECT  18.540 1.190 18.660 1.590 ;
        RECT  18.660 1.190 18.900 3.430 ;
        RECT  18.900 3.030 18.930 3.430 ;
        RECT  18.900 1.190 18.940 1.590 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.330 2.270 1.840 2.670 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  10.100 2.330 10.740 2.720 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 2.750 5.440 ;
        RECT  2.750 4.480 3.150 5.440 ;
        RECT  3.150 4.640 5.890 5.440 ;
        RECT  5.890 4.480 6.290 5.440 ;
        RECT  6.290 4.640 7.300 5.440 ;
        RECT  7.300 4.480 7.700 5.440 ;
        RECT  10.790 3.520 11.190 3.850 ;
        RECT  11.190 3.610 12.960 3.850 ;
        RECT  12.960 3.460 13.200 3.850 ;
        RECT  7.700 4.640 14.680 5.440 ;
        RECT  13.200 3.460 14.680 3.700 ;
        RECT  14.680 3.460 14.920 5.440 ;
        RECT  14.920 4.640 15.520 5.440 ;
        RECT  15.520 3.580 15.530 5.440 ;
        RECT  15.530 3.460 15.930 5.440 ;
        RECT  15.930 3.580 15.940 5.440 ;
        RECT  15.940 4.640 17.700 5.440 ;
        RECT  17.700 3.460 18.100 5.440 ;
        RECT  18.100 4.640 19.140 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.440 0.400 ;
        RECT  0.440 -0.400 0.450 0.750 ;
        RECT  0.450 -0.400 0.850 0.950 ;
        RECT  0.850 -0.400 0.860 0.750 ;
        RECT  0.860 -0.400 2.890 0.400 ;
        RECT  2.890 -0.400 3.290 0.560 ;
        RECT  3.290 -0.400 5.870 0.400 ;
        RECT  5.870 -0.400 5.880 0.730 ;
        RECT  5.880 -0.400 6.280 0.930 ;
        RECT  6.280 -0.400 6.290 0.730 ;
        RECT  6.290 -0.400 8.810 0.400 ;
        RECT  8.810 -0.400 8.820 0.730 ;
        RECT  8.820 -0.400 9.220 0.850 ;
        RECT  9.220 -0.400 9.230 0.730 ;
        RECT  9.230 -0.400 10.900 0.400 ;
        RECT  10.900 -0.400 10.910 1.420 ;
        RECT  10.910 -0.400 11.310 1.540 ;
        RECT  11.310 -0.400 11.320 1.420 ;
        RECT  11.320 -0.400 13.460 0.400 ;
        RECT  13.460 -0.400 13.860 0.560 ;
        RECT  13.860 -0.400 17.700 0.400 ;
        RECT  17.700 -0.400 17.710 0.990 ;
        RECT  17.710 -0.400 18.110 1.480 ;
        RECT  18.110 -0.400 18.120 0.990 ;
        RECT  18.120 -0.400 19.140 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  18.020 1.870 18.420 2.270 ;
        RECT  17.150 1.950 18.020 2.190 ;
        RECT  16.910 1.390 17.150 3.170 ;
        RECT  15.870 0.780 16.110 1.500 ;
        RECT  15.430 2.250 16.050 2.650 ;
        RECT  14.670 0.780 15.870 1.020 ;
        RECT  15.190 1.310 15.430 3.170 ;
        RECT  15.030 1.310 15.190 1.550 ;
        RECT  13.530 2.930 15.190 3.170 ;
        RECT  14.630 1.850 14.870 2.260 ;
        RECT  14.430 0.780 14.670 1.500 ;
        RECT  12.680 1.850 14.630 2.090 ;
        RECT  14.270 1.100 14.430 1.500 ;
        RECT  13.130 2.600 13.530 3.170 ;
        RECT  11.900 0.730 13.030 0.970 ;
        RECT  12.440 1.290 12.680 3.330 ;
        RECT  12.180 1.290 12.440 1.530 ;
        RECT  12.090 3.090 12.440 3.330 ;
        RECT  11.890 2.520 12.160 2.760 ;
        RECT  11.890 0.730 11.900 2.060 ;
        RECT  11.810 0.730 11.890 2.760 ;
        RECT  11.650 0.730 11.810 3.230 ;
        RECT  11.570 1.820 11.650 3.230 ;
        RECT  11.560 1.820 11.570 2.590 ;
        RECT  10.430 2.990 11.570 3.230 ;
        RECT  10.430 1.820 11.560 2.060 ;
        RECT  10.190 1.460 10.430 2.060 ;
        RECT  10.190 2.990 10.430 3.840 ;
        RECT  9.750 0.770 10.260 1.010 ;
        RECT  10.030 1.460 10.190 1.700 ;
        RECT  10.030 3.430 10.190 3.840 ;
        RECT  8.710 3.600 10.030 3.840 ;
        RECT  9.510 0.770 9.750 1.370 ;
        RECT  9.500 1.650 9.740 3.140 ;
        RECT  7.820 1.130 9.510 1.370 ;
        RECT  9.030 1.650 9.500 1.890 ;
        RECT  9.390 2.900 9.500 3.140 ;
        RECT  8.990 2.900 9.390 3.320 ;
        RECT  8.260 2.900 8.990 3.140 ;
        RECT  8.470 3.420 8.710 3.840 ;
        RECT  5.540 3.420 8.470 3.660 ;
        RECT  8.020 2.510 8.260 3.140 ;
        RECT  7.740 1.090 7.820 1.490 ;
        RECT  7.500 1.090 7.740 3.140 ;
        RECT  7.420 1.090 7.500 1.490 ;
        RECT  6.060 2.900 7.500 3.140 ;
        RECT  6.980 1.780 7.220 2.180 ;
        RECT  5.490 1.940 6.980 2.180 ;
        RECT  5.820 2.460 6.060 3.140 ;
        RECT  5.300 3.420 5.540 4.360 ;
        RECT  5.250 1.070 5.490 2.680 ;
        RECT  5.050 4.120 5.300 4.360 ;
        RECT  5.240 1.070 5.250 2.180 ;
        RECT  4.990 2.440 5.250 2.680 ;
        RECT  4.910 1.070 5.240 1.310 ;
        RECT  4.990 3.450 5.020 3.850 ;
        RECT  4.780 2.440 4.990 3.850 ;
        RECT  4.720 1.740 4.960 2.140 ;
        RECT  4.510 0.910 4.910 1.310 ;
        RECT  4.750 2.440 4.780 3.840 ;
        RECT  4.370 1.740 4.720 1.980 ;
        RECT  4.370 3.250 4.450 3.650 ;
        RECT  4.130 1.740 4.370 3.650 ;
        RECT  4.030 1.740 4.130 1.980 ;
        RECT  3.560 3.300 4.130 3.650 ;
        RECT  3.630 0.660 4.030 1.100 ;
        RECT  3.630 1.410 4.030 1.980 ;
        RECT  3.940 3.970 4.020 4.370 ;
        RECT  3.620 3.940 3.940 4.370 ;
        RECT  2.260 0.860 3.630 1.100 ;
        RECT  3.260 3.940 3.620 4.180 ;
        RECT  3.020 3.610 3.260 4.180 ;
        RECT  2.020 3.610 3.020 3.850 ;
        RECT  2.020 0.860 2.260 1.590 ;
        RECT  1.090 4.130 2.180 4.370 ;
        RECT  1.950 1.350 2.020 1.590 ;
        RECT  1.780 3.340 2.020 3.850 ;
        RECT  1.710 1.350 1.950 1.750 ;
        RECT  1.620 3.340 1.780 3.580 ;
        RECT  1.360 0.670 1.730 0.910 ;
        RECT  1.120 0.670 1.360 1.990 ;
        RECT  0.930 1.750 1.120 1.990 ;
        RECT  0.850 3.940 1.090 4.370 ;
        RECT  0.690 1.750 0.930 2.360 ;
        RECT  0.400 3.940 0.850 4.180 ;
        RECT  0.400 2.120 0.690 2.360 ;
        RECT  0.160 2.120 0.400 4.180 ;
    END
END SDFFSRX1

MACRO SDFFSHQXL
    CLASS CORE ;
    FOREIGN SDFFSHQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.970 2.530 7.210 2.930 ;
        RECT  7.210 2.530 7.460 2.860 ;
        RECT  7.460 2.390 7.720 2.860 ;
        RECT  7.720 2.620 7.940 2.860 ;
        RECT  7.940 2.620 8.180 4.180 ;
        RECT  8.180 3.940 9.800 4.180 ;
        RECT  9.800 3.940 10.040 4.370 ;
        RECT  10.040 4.080 10.110 4.370 ;
        RECT  10.110 4.130 13.650 4.370 ;
        RECT  13.650 4.080 13.790 4.370 ;
        RECT  13.790 2.160 13.930 4.370 ;
        RECT  13.930 2.080 14.030 4.370 ;
        RECT  14.030 2.080 14.070 2.640 ;
        RECT  14.070 2.080 14.330 2.480 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.770 2.360 2.780 2.650 ;
        RECT  2.780 2.190 3.180 2.650 ;
        RECT  3.180 2.360 3.190 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.410 2.380 1.870 2.810 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.470 3.220 14.630 3.620 ;
        RECT  14.630 2.790 14.870 3.620 ;
        RECT  14.870 2.790 15.290 3.030 ;
        RECT  15.290 2.660 15.390 3.030 ;
        RECT  15.380 1.830 15.390 2.090 ;
        RECT  15.350 1.000 15.390 1.400 ;
        RECT  15.390 1.000 15.630 3.030 ;
        RECT  15.630 1.830 15.640 2.090 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.980 1.740 4.510 2.160 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.040 0.780 2.440 ;
        RECT  0.780 1.840 0.860 2.440 ;
        RECT  0.860 1.830 1.030 2.440 ;
        RECT  1.030 1.830 1.120 2.090 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.200 5.440 ;
        RECT  0.200 4.480 0.600 5.440 ;
        RECT  0.600 4.640 3.700 5.440 ;
        RECT  3.700 4.110 3.940 5.440 ;
        RECT  3.940 4.640 6.690 5.440 ;
        RECT  6.690 4.090 7.670 5.440 ;
        RECT  7.670 4.640 9.110 5.440 ;
        RECT  9.110 4.480 9.510 5.440 ;
        RECT  9.510 4.640 14.310 5.440 ;
        RECT  14.310 4.480 14.710 5.440 ;
        RECT  14.710 4.640 15.220 5.440 ;
        RECT  15.220 3.510 15.230 5.440 ;
        RECT  15.230 3.310 15.630 5.440 ;
        RECT  15.630 3.510 15.640 5.440 ;
        RECT  15.640 4.640 15.840 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.830 0.400 ;
        RECT  0.830 -0.400 1.230 0.560 ;
        RECT  1.230 -0.400 2.910 0.400 ;
        RECT  2.910 -0.400 3.310 0.560 ;
        RECT  3.310 -0.400 6.340 0.400 ;
        RECT  6.340 -0.400 6.350 0.730 ;
        RECT  6.350 -0.400 6.750 0.850 ;
        RECT  6.750 -0.400 6.760 0.730 ;
        RECT  6.760 -0.400 9.390 0.400 ;
        RECT  9.390 -0.400 9.630 1.300 ;
        RECT  9.630 -0.400 12.350 0.400 ;
        RECT  12.350 -0.400 12.750 0.560 ;
        RECT  12.750 -0.400 13.990 0.400 ;
        RECT  13.990 -0.400 14.390 0.560 ;
        RECT  14.390 -0.400 15.840 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.770 1.280 15.010 2.510 ;
        RECT  13.770 1.280 14.770 1.520 ;
        RECT  13.530 0.860 13.770 1.520 ;
        RECT  13.430 0.860 13.530 1.100 ;
        RECT  12.610 3.590 13.450 3.830 ;
        RECT  13.030 0.690 13.430 1.100 ;
        RECT  12.510 0.860 13.030 1.100 ;
        RECT  12.790 1.380 13.030 2.710 ;
        RECT  12.610 2.470 12.790 2.710 ;
        RECT  12.370 2.470 12.610 3.830 ;
        RECT  12.270 0.860 12.510 2.190 ;
        RECT  12.070 0.860 12.270 1.100 ;
        RECT  12.090 1.950 12.270 2.190 ;
        RECT  11.850 1.950 12.090 3.130 ;
        RECT  11.780 0.780 12.070 1.100 ;
        RECT  10.860 2.890 11.850 3.130 ;
        RECT  9.450 3.410 11.830 3.650 ;
        RECT  11.010 0.780 11.780 1.020 ;
        RECT  11.440 1.380 11.730 1.620 ;
        RECT  11.200 1.380 11.440 2.370 ;
        RECT  10.490 2.130 11.200 2.370 ;
        RECT  10.430 1.010 10.590 1.410 ;
        RECT  10.250 2.130 10.490 2.610 ;
        RECT  10.190 1.010 10.430 1.840 ;
        RECT  9.970 2.890 10.380 3.130 ;
        RECT  9.970 1.600 10.190 1.840 ;
        RECT  9.730 1.600 9.970 3.130 ;
        RECT  9.210 1.580 9.450 3.650 ;
        RECT  9.110 1.580 9.210 1.820 ;
        RECT  8.510 3.410 9.210 3.650 ;
        RECT  8.870 1.350 9.110 1.820 ;
        RECT  8.680 2.110 8.920 2.690 ;
        RECT  8.750 1.350 8.870 1.590 ;
        RECT  8.510 0.670 8.750 1.590 ;
        RECT  8.590 2.110 8.680 2.350 ;
        RECT  8.350 1.870 8.590 2.350 ;
        RECT  8.290 0.670 8.510 0.910 ;
        RECT  8.090 1.870 8.350 2.110 ;
        RECT  7.850 1.350 8.090 2.110 ;
        RECT  7.690 1.350 7.850 2.080 ;
        RECT  7.410 0.770 7.790 1.010 ;
        RECT  6.690 1.840 7.690 2.080 ;
        RECT  6.690 3.370 7.470 3.610 ;
        RECT  7.170 0.770 7.410 1.370 ;
        RECT  5.930 1.130 7.170 1.370 ;
        RECT  6.450 1.840 6.690 3.610 ;
        RECT  6.170 1.840 6.450 2.080 ;
        RECT  5.930 2.360 6.170 4.050 ;
        RECT  5.890 0.940 5.930 1.370 ;
        RECT  5.890 2.360 5.930 2.600 ;
        RECT  5.190 3.810 5.930 4.050 ;
        RECT  5.650 0.940 5.890 2.600 ;
        RECT  5.010 0.940 5.650 1.180 ;
        RECT  5.410 3.040 5.650 3.440 ;
        RECT  5.190 3.040 5.410 3.280 ;
        RECT  4.950 1.880 5.190 3.280 ;
        RECT  4.010 2.710 4.950 2.950 ;
        RECT  4.370 3.230 4.610 3.830 ;
        RECT  2.630 0.890 4.590 1.130 ;
        RECT  3.420 3.590 4.370 3.830 ;
        RECT  3.770 2.710 4.010 3.310 ;
        RECT  2.900 3.070 3.770 3.310 ;
        RECT  2.380 1.470 3.620 1.710 ;
        RECT  3.180 3.590 3.420 4.370 ;
        RECT  1.770 4.130 3.180 4.370 ;
        RECT  2.660 3.070 2.900 3.850 ;
        RECT  0.580 3.610 2.660 3.850 ;
        RECT  2.390 0.670 2.630 1.130 ;
        RECT  1.570 0.670 2.390 0.910 ;
        RECT  2.140 1.470 2.380 3.320 ;
        RECT  1.710 1.470 2.140 1.870 ;
        RECT  1.650 3.080 2.140 3.320 ;
        RECT  0.400 3.080 0.580 3.850 ;
        RECT  0.400 1.360 0.490 1.760 ;
        RECT  0.340 1.360 0.400 3.850 ;
        RECT  0.160 1.360 0.340 3.320 ;
    END
END SDFFSHQXL

MACRO SDFFSHQX4
    CLASS CORE ;
    FOREIGN SDFFSHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSHQXL ;
    SIZE 21.120 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.130 2.400 7.460 2.880 ;
        RECT  7.460 2.390 7.720 2.880 ;
        RECT  7.720 2.640 8.230 2.880 ;
        RECT  8.230 2.640 8.470 3.660 ;
        RECT  8.470 3.420 10.490 3.660 ;
        RECT  10.490 3.420 10.730 3.730 ;
        RECT  10.730 3.490 12.150 3.730 ;
        RECT  12.150 3.490 12.390 4.180 ;
        RECT  12.390 3.620 12.430 4.180 ;
        RECT  12.430 3.940 17.270 4.180 ;
        RECT  17.270 3.640 17.580 4.180 ;
        RECT  17.580 2.260 17.820 4.180 ;
        RECT  17.820 2.260 18.010 2.660 ;
        RECT  18.010 2.360 19.210 2.660 ;
        RECT  19.210 2.250 19.560 2.660 ;
        RECT  19.560 2.250 19.610 2.650 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.810 2.550 2.840 2.790 ;
        RECT  2.840 2.390 2.850 2.790 ;
        RECT  2.690 1.380 2.850 1.830 ;
        RECT  2.850 1.380 3.090 2.790 ;
        RECT  3.090 2.390 3.100 2.790 ;
        RECT  3.100 2.550 3.210 2.790 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.260 2.380 1.720 2.810 ;
        RECT  1.720 2.390 1.770 2.720 ;
        RECT  1.770 2.390 1.780 2.650 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.110 0.800 18.510 1.390 ;
        RECT  18.170 3.050 18.570 4.030 ;
        RECT  18.570 3.050 18.810 3.300 ;
        RECT  18.810 3.060 19.550 3.300 ;
        RECT  19.550 2.940 19.690 3.300 ;
        RECT  19.690 2.940 19.910 4.050 ;
        RECT  19.910 2.940 20.350 4.340 ;
        RECT  18.510 1.150 20.550 1.390 ;
        RECT  20.350 2.940 20.710 3.220 ;
        RECT  20.550 0.770 20.710 1.390 ;
        RECT  20.710 0.770 20.800 3.220 ;
        RECT  20.800 0.770 20.950 3.190 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.880 1.640 4.430 2.090 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.690 1.830 0.930 2.360 ;
        RECT  0.930 1.830 1.180 2.090 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 4.480 1.390 5.440 ;
        RECT  1.390 4.640 3.700 5.440 ;
        RECT  3.700 4.110 3.940 5.440 ;
        RECT  3.940 4.640 6.720 5.440 ;
        RECT  6.720 4.480 7.120 5.440 ;
        RECT  7.120 4.640 8.360 5.440 ;
        RECT  8.360 4.480 8.760 5.440 ;
        RECT  8.760 4.640 9.790 5.440 ;
        RECT  9.790 4.060 9.800 5.440 ;
        RECT  9.800 3.940 10.200 5.440 ;
        RECT  10.200 4.060 10.210 5.440 ;
        RECT  10.210 4.640 11.440 5.440 ;
        RECT  11.440 4.130 11.450 5.440 ;
        RECT  11.450 4.010 11.850 5.440 ;
        RECT  11.850 4.130 11.860 5.440 ;
        RECT  11.860 4.640 15.890 5.440 ;
        RECT  15.890 4.480 16.290 5.440 ;
        RECT  16.290 4.640 17.350 5.440 ;
        RECT  17.350 4.480 17.750 5.440 ;
        RECT  17.750 4.640 18.920 5.440 ;
        RECT  18.920 4.090 18.930 5.440 ;
        RECT  18.930 3.600 19.330 5.440 ;
        RECT  19.330 4.090 19.340 5.440 ;
        RECT  19.340 4.640 20.620 5.440 ;
        RECT  20.620 3.600 20.860 5.440 ;
        RECT  20.860 4.640 21.120 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.920 0.400 ;
        RECT  0.920 -0.400 0.930 1.080 ;
        RECT  0.930 -0.400 1.330 1.280 ;
        RECT  1.330 -0.400 1.340 1.080 ;
        RECT  1.340 -0.400 3.010 0.400 ;
        RECT  3.010 -0.400 3.410 0.560 ;
        RECT  3.410 -0.400 6.420 0.400 ;
        RECT  6.420 -0.400 6.430 0.730 ;
        RECT  6.430 -0.400 6.830 0.850 ;
        RECT  6.830 -0.400 6.840 0.730 ;
        RECT  6.840 -0.400 9.900 0.400 ;
        RECT  9.900 -0.400 9.910 1.320 ;
        RECT  9.910 -0.400 10.310 1.440 ;
        RECT  10.310 -0.400 10.320 1.320 ;
        RECT  10.320 -0.400 11.420 0.400 ;
        RECT  11.420 -0.400 11.430 1.110 ;
        RECT  11.430 -0.400 11.830 1.230 ;
        RECT  11.830 -0.400 11.840 1.110 ;
        RECT  11.840 -0.400 15.660 0.400 ;
        RECT  15.660 -0.400 16.060 0.560 ;
        RECT  16.060 -0.400 16.830 0.400 ;
        RECT  16.830 -0.400 17.230 0.560 ;
        RECT  17.230 -0.400 19.320 0.400 ;
        RECT  19.320 -0.400 19.330 0.660 ;
        RECT  19.330 -0.400 19.730 0.860 ;
        RECT  19.730 -0.400 19.740 0.660 ;
        RECT  19.740 -0.400 21.120 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  20.270 2.070 20.430 2.470 ;
        RECT  20.030 1.730 20.270 2.470 ;
        RECT  17.660 1.730 20.030 1.970 ;
        RECT  17.420 0.860 17.660 1.970 ;
        RECT  14.880 0.860 17.420 1.100 ;
        RECT  16.850 1.540 17.090 3.290 ;
        RECT  16.180 1.540 16.850 1.780 ;
        RECT  16.690 2.890 16.850 3.290 ;
        RECT  16.350 2.220 16.510 2.620 ;
        RECT  16.110 2.220 16.350 3.660 ;
        RECT  15.980 1.380 16.180 1.780 ;
        RECT  14.870 3.420 16.110 3.660 ;
        RECT  15.770 1.370 15.980 1.790 ;
        RECT  15.760 1.370 15.770 2.150 ;
        RECT  15.360 1.370 15.760 2.350 ;
        RECT  15.350 1.370 15.360 2.150 ;
        RECT  14.870 0.860 14.880 1.630 ;
        RECT  14.720 0.860 14.870 3.660 ;
        RECT  14.630 0.670 14.720 3.660 ;
        RECT  14.480 0.670 14.630 1.630 ;
        RECT  13.030 3.420 14.630 3.660 ;
        RECT  13.360 0.670 14.480 0.910 ;
        RECT  13.390 2.900 14.190 3.140 ;
        RECT  13.720 1.250 14.120 1.750 ;
        RECT  13.390 1.510 13.720 1.750 ;
        RECT  13.150 1.510 13.390 3.140 ;
        RECT  13.120 0.670 13.360 1.220 ;
        RECT  12.600 1.510 13.150 1.750 ;
        RECT  12.670 2.900 13.150 3.140 ;
        RECT  12.960 0.980 13.120 1.220 ;
        RECT  10.310 2.030 12.870 2.270 ;
        RECT  12.270 2.900 12.670 3.210 ;
        RECT  12.590 1.410 12.600 1.750 ;
        RECT  12.190 1.070 12.590 1.750 ;
        RECT  10.630 2.900 12.270 3.140 ;
        RECT  11.070 1.510 12.190 1.750 ;
        RECT  10.750 1.070 11.070 1.750 ;
        RECT  10.670 1.070 10.750 1.470 ;
        RECT  10.070 1.800 10.310 3.140 ;
        RECT  9.580 1.800 10.070 2.040 ;
        RECT  9.240 2.900 10.070 3.140 ;
        RECT  8.990 2.320 9.790 2.560 ;
        RECT  9.470 1.270 9.580 2.040 ;
        RECT  9.340 0.670 9.470 2.040 ;
        RECT  9.040 3.940 9.440 4.370 ;
        RECT  9.230 0.670 9.340 1.590 ;
        RECT  8.820 0.670 9.230 0.910 ;
        RECT  6.310 3.940 9.040 4.180 ;
        RECT  8.750 1.870 8.990 2.560 ;
        RECT  8.170 1.870 8.750 2.110 ;
        RECT  7.430 0.770 8.500 1.010 ;
        RECT  7.930 1.460 8.170 2.110 ;
        RECT  6.840 3.190 7.940 3.430 ;
        RECT  7.770 1.460 7.930 1.890 ;
        RECT  6.840 1.650 7.770 1.890 ;
        RECT  7.190 0.770 7.430 1.370 ;
        RECT  5.910 1.130 7.190 1.370 ;
        RECT  6.600 1.650 6.840 3.430 ;
        RECT  6.440 1.650 6.600 2.060 ;
        RECT  6.190 1.650 6.440 2.050 ;
        RECT  5.990 3.700 6.310 4.180 ;
        RECT  5.390 3.700 5.990 3.940 ;
        RECT  5.670 0.730 5.910 3.290 ;
        RECT  5.050 0.730 5.670 0.970 ;
        RECT  5.150 2.370 5.390 3.940 ;
        RECT  5.070 2.370 5.150 2.610 ;
        RECT  4.830 1.380 5.070 2.610 ;
        RECT  4.630 2.890 4.870 3.830 ;
        RECT  3.870 2.370 4.830 2.610 ;
        RECT  3.930 0.740 4.690 0.980 ;
        RECT  3.420 3.590 4.630 3.830 ;
        RECT  3.690 0.740 3.930 1.100 ;
        RECT  3.630 2.370 3.870 3.310 ;
        RECT  2.730 0.860 3.690 1.100 ;
        RECT  2.900 3.070 3.630 3.310 ;
        RECT  3.180 3.590 3.420 4.370 ;
        RECT  1.930 4.130 3.180 4.370 ;
        RECT  2.660 3.070 2.900 3.840 ;
        RECT  2.490 0.670 2.730 1.100 ;
        RECT  0.570 3.600 2.660 3.840 ;
        RECT  1.670 0.670 2.490 0.910 ;
        RECT  2.140 1.470 2.380 3.320 ;
        RECT  1.810 1.470 2.140 1.870 ;
        RECT  1.810 3.080 2.140 3.320 ;
        RECT  0.410 1.150 0.570 1.550 ;
        RECT  0.410 2.980 0.570 3.960 ;
        RECT  0.170 1.150 0.410 3.960 ;
    END
END SDFFSHQX4

MACRO SDFFSHQX2
    CLASS CORE ;
    FOREIGN SDFFSHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSHQXL ;
    SIZE 17.820 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.970 2.400 7.210 2.810 ;
        RECT  7.210 2.400 7.460 2.690 ;
        RECT  7.460 2.390 7.720 2.690 ;
        RECT  7.720 2.450 7.750 2.690 ;
        RECT  7.750 2.450 7.940 3.110 ;
        RECT  7.940 2.450 7.990 4.360 ;
        RECT  7.990 2.870 8.180 4.360 ;
        RECT  8.180 4.120 9.690 4.360 ;
        RECT  9.690 4.080 9.770 4.360 ;
        RECT  9.770 3.650 10.010 4.360 ;
        RECT  10.010 3.650 11.050 3.890 ;
        RECT  11.050 3.650 11.290 4.370 ;
        RECT  11.290 4.060 11.430 4.370 ;
        RECT  11.430 4.130 15.450 4.370 ;
        RECT  15.450 2.270 15.690 4.370 ;
        RECT  15.690 2.270 15.850 2.670 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.820 2.300 3.340 2.760 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.340 1.820 1.780 2.270 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.250 1.390 17.370 1.790 ;
        RECT  16.580 2.880 17.410 3.280 ;
        RECT  17.370 1.390 17.410 1.840 ;
        RECT  17.410 1.390 17.650 3.280 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.120 1.670 4.540 2.230 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.340 0.770 2.740 ;
        RECT  0.770 2.340 0.860 3.200 ;
        RECT  0.860 2.340 1.020 3.210 ;
        RECT  1.020 2.950 1.120 3.210 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.280 5.440 ;
        RECT  0.280 4.480 0.680 5.440 ;
        RECT  0.680 4.640 3.330 5.440 ;
        RECT  3.330 4.110 3.570 5.440 ;
        RECT  3.570 4.640 6.690 5.440 ;
        RECT  6.690 4.110 7.670 5.440 ;
        RECT  7.670 4.640 10.340 5.440 ;
        RECT  10.340 4.170 10.740 5.440 ;
        RECT  10.740 4.640 15.960 5.440 ;
        RECT  15.960 4.360 15.970 5.440 ;
        RECT  15.970 4.160 16.370 5.440 ;
        RECT  16.370 4.360 16.380 5.440 ;
        RECT  16.380 4.640 17.200 5.440 ;
        RECT  17.200 4.340 17.210 5.440 ;
        RECT  17.210 4.140 17.610 5.440 ;
        RECT  17.610 4.340 17.620 5.440 ;
        RECT  17.620 4.640 17.820 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.320 0.400 ;
        RECT  0.320 -0.400 0.720 0.560 ;
        RECT  0.720 -0.400 2.910 0.400 ;
        RECT  2.910 -0.400 3.310 0.560 ;
        RECT  3.310 -0.400 6.320 0.400 ;
        RECT  6.320 -0.400 6.330 0.730 ;
        RECT  6.330 -0.400 6.730 0.850 ;
        RECT  6.730 -0.400 6.740 0.730 ;
        RECT  6.740 -0.400 9.310 0.400 ;
        RECT  9.310 -0.400 9.550 1.310 ;
        RECT  9.550 -0.400 10.740 0.400 ;
        RECT  10.740 -0.400 10.750 1.110 ;
        RECT  10.750 -0.400 11.150 1.310 ;
        RECT  11.150 -0.400 11.160 1.110 ;
        RECT  11.160 -0.400 14.350 0.400 ;
        RECT  14.350 -0.400 14.750 0.560 ;
        RECT  14.750 -0.400 15.980 0.400 ;
        RECT  15.980 -0.400 16.380 0.560 ;
        RECT  16.380 -0.400 17.820 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.890 2.070 17.130 2.470 ;
        RECT  16.740 2.070 16.890 2.310 ;
        RECT  16.500 0.860 16.740 2.310 ;
        RECT  13.710 0.860 16.500 1.100 ;
        RECT  14.820 2.120 15.010 3.850 ;
        RECT  14.810 1.790 14.820 3.850 ;
        RECT  14.770 1.390 14.810 3.850 ;
        RECT  14.450 1.390 14.770 2.360 ;
        RECT  14.510 3.610 14.770 3.850 ;
        RECT  13.710 2.810 14.490 3.050 ;
        RECT  14.410 1.390 14.450 2.410 ;
        RECT  14.400 1.790 14.410 2.410 ;
        RECT  14.050 2.010 14.400 2.410 ;
        RECT  13.500 0.860 13.710 3.850 ;
        RECT  13.470 0.850 13.500 3.850 ;
        RECT  13.250 0.850 13.470 1.640 ;
        RECT  11.910 3.610 13.470 3.850 ;
        RECT  13.170 0.790 13.250 1.640 ;
        RECT  12.680 3.090 13.190 3.330 ;
        RECT  13.010 0.790 13.170 1.630 ;
        RECT  11.890 0.790 13.010 1.030 ;
        RECT  12.440 1.310 12.680 3.330 ;
        RECT  12.210 1.310 12.440 1.830 ;
        RECT  11.550 3.090 12.440 3.330 ;
        RECT  10.390 1.590 12.210 1.830 ;
        RECT  9.450 2.110 12.130 2.350 ;
        RECT  11.490 0.790 11.890 1.310 ;
        RECT  11.230 3.090 11.550 3.370 ;
        RECT  9.730 3.130 11.230 3.370 ;
        RECT  10.150 0.910 10.390 1.830 ;
        RECT  9.990 0.910 10.150 1.310 ;
        RECT  9.210 1.590 9.450 3.840 ;
        RECT  9.030 1.590 9.210 1.830 ;
        RECT  8.510 3.360 9.210 3.760 ;
        RECT  8.790 1.350 9.030 1.830 ;
        RECT  8.690 2.110 8.930 2.610 ;
        RECT  8.670 1.350 8.790 1.590 ;
        RECT  8.510 2.110 8.690 2.350 ;
        RECT  8.430 0.670 8.670 1.590 ;
        RECT  8.270 1.870 8.510 2.350 ;
        RECT  8.210 0.670 8.430 0.910 ;
        RECT  8.010 1.870 8.270 2.110 ;
        RECT  7.770 1.350 8.010 2.110 ;
        RECT  7.250 0.770 7.770 1.010 ;
        RECT  7.720 1.350 7.770 1.900 ;
        RECT  7.610 1.350 7.720 1.890 ;
        RECT  6.670 1.650 7.610 1.890 ;
        RECT  7.070 3.210 7.470 3.610 ;
        RECT  7.010 0.770 7.250 1.370 ;
        RECT  6.670 3.290 7.070 3.530 ;
        RECT  5.620 1.130 7.010 1.370 ;
        RECT  6.430 1.650 6.670 3.530 ;
        RECT  6.090 2.140 6.430 2.540 ;
        RECT  4.990 4.060 5.830 4.300 ;
        RECT  5.380 0.670 5.620 3.600 ;
        RECT  4.990 0.670 5.380 0.910 ;
        RECT  5.270 3.200 5.380 3.600 ;
        RECT  4.990 1.820 5.100 2.910 ;
        RECT  4.860 1.820 4.990 4.300 ;
        RECT  4.750 2.670 4.860 4.300 ;
        RECT  2.530 3.070 4.750 3.310 ;
        RECT  4.490 0.670 4.650 0.910 ;
        RECT  4.250 0.670 4.490 1.100 ;
        RECT  4.230 3.590 4.470 4.090 ;
        RECT  2.630 0.860 4.250 1.100 ;
        RECT  3.050 3.590 4.230 3.830 ;
        RECT  2.470 1.670 3.740 1.910 ;
        RECT  2.810 3.590 3.050 4.360 ;
        RECT  1.770 4.120 2.810 4.360 ;
        RECT  2.390 0.670 2.630 1.100 ;
        RECT  2.290 3.070 2.530 3.840 ;
        RECT  2.380 1.670 2.470 2.790 ;
        RECT  1.570 0.670 2.390 0.910 ;
        RECT  2.230 1.450 2.380 2.790 ;
        RECT  0.490 3.600 2.290 3.840 ;
        RECT  2.140 1.450 2.230 1.910 ;
        RECT  1.970 2.550 2.230 2.790 ;
        RECT  1.730 2.550 1.970 3.320 ;
        RECT  0.400 1.250 0.490 1.650 ;
        RECT  0.400 3.080 0.490 3.840 ;
        RECT  0.250 1.250 0.400 3.840 ;
        RECT  0.160 1.250 0.250 3.400 ;
    END
END SDFFSHQX2

MACRO SDFFSHQX1
    CLASS CORE ;
    FOREIGN SDFFSHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSHQXL ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.970 2.550 7.460 2.950 ;
        RECT  7.460 2.390 7.720 2.950 ;
        RECT  7.720 2.660 7.940 2.950 ;
        RECT  7.940 2.660 8.180 4.180 ;
        RECT  8.180 3.940 9.800 4.180 ;
        RECT  9.800 3.930 10.110 4.180 ;
        RECT  10.110 3.930 13.930 4.170 ;
        RECT  13.930 2.080 14.170 4.170 ;
        RECT  14.170 2.080 14.330 2.480 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.660 1.380 2.750 1.620 ;
        RECT  2.810 2.540 2.840 2.780 ;
        RECT  2.840 2.390 2.850 2.780 ;
        RECT  2.750 1.380 2.850 1.820 ;
        RECT  2.850 1.380 3.090 2.780 ;
        RECT  3.090 2.390 3.100 2.780 ;
        RECT  3.100 2.540 3.210 2.780 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.410 2.380 1.870 2.810 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.470 3.070 14.690 3.470 ;
        RECT  14.690 2.820 14.930 3.470 ;
        RECT  14.930 2.820 15.290 3.060 ;
        RECT  15.290 2.620 15.390 3.060 ;
        RECT  15.380 1.830 15.390 2.090 ;
        RECT  15.270 0.870 15.390 1.270 ;
        RECT  15.390 0.870 15.630 3.060 ;
        RECT  15.630 2.620 15.640 2.870 ;
        RECT  15.630 1.830 15.640 2.090 ;
        RECT  15.630 0.870 15.670 1.390 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.890 1.770 4.420 2.250 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.040 0.780 2.540 ;
        RECT  0.780 1.840 0.860 2.540 ;
        RECT  0.860 1.830 0.920 2.540 ;
        RECT  0.920 1.830 1.020 2.280 ;
        RECT  1.020 1.830 1.120 2.090 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.780 5.440 ;
        RECT  0.780 4.480 1.180 5.440 ;
        RECT  1.180 4.640 3.700 5.440 ;
        RECT  3.700 4.110 3.940 5.440 ;
        RECT  3.940 4.640 6.630 5.440 ;
        RECT  6.630 4.110 7.610 5.440 ;
        RECT  7.610 4.640 9.110 5.440 ;
        RECT  9.110 4.480 9.510 5.440 ;
        RECT  9.510 4.640 12.520 5.440 ;
        RECT  12.520 4.480 14.060 5.440 ;
        RECT  14.060 4.640 15.220 5.440 ;
        RECT  15.220 3.540 15.230 5.440 ;
        RECT  15.230 3.340 15.630 5.440 ;
        RECT  15.630 3.540 15.640 5.440 ;
        RECT  15.640 4.640 15.840 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.760 0.400 ;
        RECT  0.760 -0.400 0.770 0.760 ;
        RECT  0.770 -0.400 1.170 0.960 ;
        RECT  1.170 -0.400 1.180 0.760 ;
        RECT  1.180 -0.400 2.850 0.400 ;
        RECT  2.850 -0.400 3.250 0.560 ;
        RECT  3.250 -0.400 6.340 0.400 ;
        RECT  6.340 -0.400 6.350 0.730 ;
        RECT  6.350 -0.400 6.750 0.850 ;
        RECT  6.750 -0.400 6.760 0.730 ;
        RECT  6.760 -0.400 9.390 0.400 ;
        RECT  9.390 -0.400 9.630 1.310 ;
        RECT  9.630 -0.400 12.330 0.400 ;
        RECT  12.330 -0.400 12.730 0.560 ;
        RECT  12.730 -0.400 14.040 0.400 ;
        RECT  14.040 -0.400 14.050 1.070 ;
        RECT  14.050 -0.400 14.450 1.270 ;
        RECT  14.450 -0.400 14.460 1.070 ;
        RECT  14.460 -0.400 15.840 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.780 1.550 15.020 2.540 ;
        RECT  13.250 1.550 14.780 1.790 ;
        RECT  13.070 2.900 13.470 3.300 ;
        RECT  13.010 0.860 13.250 2.350 ;
        RECT  12.730 2.900 13.070 3.140 ;
        RECT  12.210 0.860 13.010 1.100 ;
        RECT  12.490 1.380 12.730 3.140 ;
        RECT  11.980 2.470 12.490 2.870 ;
        RECT  12.050 0.860 12.210 2.190 ;
        RECT  11.970 0.780 12.050 2.190 ;
        RECT  10.990 0.780 11.970 1.100 ;
        RECT  11.530 1.950 11.970 2.190 ;
        RECT  11.010 1.380 11.690 1.620 ;
        RECT  9.370 3.410 11.660 3.650 ;
        RECT  11.290 1.950 11.530 3.130 ;
        RECT  10.690 2.890 11.290 3.130 ;
        RECT  10.770 1.380 11.010 2.450 ;
        RECT  10.450 2.210 10.770 2.450 ;
        RECT  10.310 1.050 10.470 1.450 ;
        RECT  10.210 2.210 10.450 2.610 ;
        RECT  9.890 2.890 10.330 3.130 ;
        RECT  10.070 1.050 10.310 1.840 ;
        RECT  9.890 1.600 10.070 1.840 ;
        RECT  9.650 1.600 9.890 3.130 ;
        RECT  9.130 1.590 9.370 3.650 ;
        RECT  9.110 1.590 9.130 1.830 ;
        RECT  9.010 3.390 9.130 3.650 ;
        RECT  8.870 1.350 9.110 1.830 ;
        RECT  8.510 3.390 9.010 3.630 ;
        RECT  8.750 1.350 8.870 1.590 ;
        RECT  8.610 2.110 8.850 2.670 ;
        RECT  8.510 0.670 8.750 1.590 ;
        RECT  8.590 2.110 8.610 2.350 ;
        RECT  8.350 1.870 8.590 2.350 ;
        RECT  8.110 0.670 8.510 0.910 ;
        RECT  8.100 1.870 8.350 2.110 ;
        RECT  7.860 1.350 8.100 2.110 ;
        RECT  7.690 1.350 7.860 2.000 ;
        RECT  7.270 0.770 7.790 1.010 ;
        RECT  6.690 1.760 7.690 2.000 ;
        RECT  6.690 3.390 7.470 3.630 ;
        RECT  7.030 0.770 7.270 1.370 ;
        RECT  5.930 1.130 7.030 1.370 ;
        RECT  6.450 1.760 6.690 3.630 ;
        RECT  6.210 1.760 6.450 2.160 ;
        RECT  5.930 2.440 6.170 4.040 ;
        RECT  5.920 0.670 5.930 1.370 ;
        RECT  5.920 2.440 5.930 2.680 ;
        RECT  5.190 3.800 5.930 4.040 ;
        RECT  5.680 0.670 5.920 2.680 ;
        RECT  4.930 0.670 5.680 0.910 ;
        RECT  5.410 2.960 5.650 3.530 ;
        RECT  5.400 2.960 5.410 3.200 ;
        RECT  5.160 2.790 5.400 3.200 ;
        RECT  5.090 2.790 5.160 3.030 ;
        RECT  4.850 1.810 5.090 3.030 ;
        RECT  4.010 2.790 4.850 3.030 ;
        RECT  4.530 3.310 4.690 3.550 ;
        RECT  4.190 0.860 4.590 1.290 ;
        RECT  4.290 3.310 4.530 3.830 ;
        RECT  3.420 3.590 4.290 3.830 ;
        RECT  1.910 0.860 4.190 1.100 ;
        RECT  3.770 2.790 4.010 3.310 ;
        RECT  2.900 3.070 3.770 3.310 ;
        RECT  3.180 3.590 3.420 4.370 ;
        RECT  1.770 4.130 3.180 4.370 ;
        RECT  2.660 3.070 2.900 3.850 ;
        RECT  0.570 3.610 2.660 3.850 ;
        RECT  2.150 1.630 2.380 3.320 ;
        RECT  2.140 1.470 2.150 3.320 ;
        RECT  1.980 1.470 2.140 1.880 ;
        RECT  1.650 3.080 2.140 3.320 ;
        RECT  1.650 1.470 1.980 1.870 ;
        RECT  1.510 0.670 1.910 1.100 ;
        RECT  0.400 3.070 0.570 3.850 ;
        RECT  0.400 1.360 0.490 1.760 ;
        RECT  0.330 1.360 0.400 3.850 ;
        RECT  0.250 1.360 0.330 3.470 ;
        RECT  0.160 1.440 0.250 3.470 ;
    END
END SDFFSHQX1

MACRO SDFFSXL
    CLASS CORE ;
    FOREIGN SDFFSXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  12.630 3.960 13.260 4.360 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.260 2.080 3.270 2.650 ;
        RECT  3.270 2.020 3.670 2.650 ;
        RECT  3.670 2.080 3.680 2.650 ;
        RECT  3.680 2.390 3.760 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.470 1.680 1.870 2.280 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.470 3.520 14.720 3.950 ;
        RECT  14.720 3.510 14.870 3.950 ;
        RECT  14.530 0.690 14.930 1.100 ;
        RECT  14.870 3.510 14.980 3.770 ;
        RECT  14.930 0.860 15.290 1.100 ;
        RECT  14.980 3.520 15.430 3.760 ;
        RECT  15.290 0.860 15.430 1.280 ;
        RECT  15.430 0.860 15.670 3.760 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.950 3.160 16.000 3.560 ;
        RECT  16.000 1.280 16.300 3.570 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.120 1.520 4.130 2.090 ;
        RECT  4.130 1.400 4.530 2.090 ;
        RECT  4.530 1.520 4.540 2.090 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.260 0.800 2.660 ;
        RECT  0.800 2.250 1.130 2.670 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.270 5.440 ;
        RECT  0.270 4.480 0.670 5.440 ;
        RECT  0.670 4.640 3.430 5.440 ;
        RECT  3.430 4.110 3.670 5.440 ;
        RECT  3.670 4.640 6.800 5.440 ;
        RECT  6.800 4.480 7.200 5.440 ;
        RECT  7.200 4.640 8.320 5.440 ;
        RECT  8.320 4.310 8.330 5.440 ;
        RECT  8.330 4.190 8.730 5.440 ;
        RECT  8.730 4.310 8.740 5.440 ;
        RECT  8.740 4.640 9.640 5.440 ;
        RECT  9.640 4.310 9.650 5.440 ;
        RECT  9.650 4.190 10.050 5.440 ;
        RECT  10.050 4.310 10.060 5.440 ;
        RECT  10.060 4.640 11.940 5.440 ;
        RECT  11.940 4.210 11.950 5.440 ;
        RECT  11.950 4.010 12.350 5.440 ;
        RECT  12.350 4.210 12.360 5.440 ;
        RECT  12.360 4.640 13.700 5.440 ;
        RECT  13.700 3.930 13.710 5.440 ;
        RECT  13.710 3.730 14.110 5.440 ;
        RECT  14.110 3.930 14.120 5.440 ;
        RECT  14.120 4.640 15.260 5.440 ;
        RECT  15.260 4.480 15.660 5.440 ;
        RECT  15.660 4.640 16.500 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.020 0.400 ;
        RECT  1.020 -0.400 1.420 0.560 ;
        RECT  1.420 -0.400 3.090 0.400 ;
        RECT  3.090 -0.400 3.490 0.560 ;
        RECT  3.490 -0.400 6.640 0.400 ;
        RECT  6.640 -0.400 6.650 0.750 ;
        RECT  6.650 -0.400 7.050 0.870 ;
        RECT  7.050 -0.400 7.060 0.750 ;
        RECT  7.060 -0.400 9.300 0.400 ;
        RECT  9.300 -0.400 9.310 0.730 ;
        RECT  9.310 -0.400 9.710 0.850 ;
        RECT  9.710 -0.400 9.720 0.730 ;
        RECT  9.720 -0.400 11.890 0.400 ;
        RECT  11.890 -0.400 12.290 0.560 ;
        RECT  12.290 -0.400 13.640 0.400 ;
        RECT  13.640 -0.400 13.650 0.850 ;
        RECT  13.650 -0.400 14.050 1.050 ;
        RECT  14.050 -0.400 14.060 0.850 ;
        RECT  14.060 -0.400 15.270 0.400 ;
        RECT  15.270 -0.400 15.670 0.560 ;
        RECT  15.670 -0.400 16.500 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.940 1.960 15.150 2.370 ;
        RECT  14.930 1.500 14.940 2.370 ;
        RECT  14.690 1.380 14.930 3.210 ;
        RECT  14.680 1.380 14.690 2.110 ;
        RECT  14.530 2.810 14.690 3.210 ;
        RECT  14.530 1.380 14.680 1.780 ;
        RECT  14.090 2.020 14.250 2.420 ;
        RECT  13.850 1.570 14.090 3.210 ;
        RECT  12.710 1.570 13.850 1.810 ;
        RECT  13.230 2.970 13.850 3.210 ;
        RECT  12.830 2.970 13.230 3.370 ;
        RECT  12.530 2.290 12.930 2.690 ;
        RECT  12.310 1.220 12.710 1.810 ;
        RECT  11.530 2.370 12.530 2.610 ;
        RECT  12.050 1.570 12.310 1.810 ;
        RECT  11.810 1.570 12.050 1.970 ;
        RECT  11.290 1.490 11.530 4.370 ;
        RECT  10.770 1.490 11.290 1.730 ;
        RECT  10.770 2.730 11.010 3.910 ;
        RECT  10.530 1.330 10.770 1.730 ;
        RECT  9.250 3.670 10.770 3.910 ;
        RECT  10.250 2.010 10.550 2.410 ;
        RECT  10.010 1.240 10.250 3.390 ;
        RECT  8.870 1.240 10.010 1.480 ;
        RECT  9.210 3.150 10.010 3.390 ;
        RECT  9.490 2.020 9.730 2.420 ;
        RECT  8.820 2.100 9.490 2.340 ;
        RECT  9.010 3.670 9.250 4.070 ;
        RECT  6.510 3.670 9.010 3.910 ;
        RECT  8.630 0.670 8.870 1.480 ;
        RECT  8.580 1.760 8.820 3.400 ;
        RECT  7.330 0.670 8.630 0.910 ;
        RECT  8.350 1.760 8.580 2.000 ;
        RECT  6.870 3.160 8.580 3.400 ;
        RECT  8.110 1.430 8.350 2.000 ;
        RECT  8.050 2.370 8.290 2.770 ;
        RECT  7.580 2.370 8.050 2.610 ;
        RECT  7.340 1.460 7.580 2.610 ;
        RECT  5.990 1.460 7.340 1.700 ;
        RECT  6.630 2.160 6.870 3.400 ;
        RECT  6.270 3.670 6.510 4.140 ;
        RECT  5.470 3.900 6.270 4.140 ;
        RECT  5.750 1.150 5.990 3.500 ;
        RECT  5.710 1.150 5.750 1.390 ;
        RECT  5.310 0.760 5.710 1.390 ;
        RECT  5.230 1.670 5.470 4.140 ;
        RECT  5.090 1.670 5.230 2.070 ;
        RECT  4.190 3.900 5.230 4.140 ;
        RECT  4.710 3.070 4.950 3.500 ;
        RECT  4.430 0.700 4.830 1.100 ;
        RECT  2.630 3.070 4.710 3.310 ;
        RECT  2.570 0.860 4.430 1.100 ;
        RECT  3.950 3.590 4.190 4.140 ;
        RECT  3.150 3.590 3.950 3.830 ;
        RECT  2.850 1.380 3.790 1.620 ;
        RECT  2.910 3.590 3.150 4.370 ;
        RECT  2.850 2.550 2.930 2.790 ;
        RECT  1.940 4.130 2.910 4.370 ;
        RECT  2.610 1.380 2.850 2.790 ;
        RECT  2.390 3.070 2.630 3.850 ;
        RECT  2.260 1.420 2.610 1.830 ;
        RECT  2.110 2.550 2.610 2.790 ;
        RECT  2.330 0.670 2.570 1.100 ;
        RECT  2.230 3.610 2.390 3.850 ;
        RECT  1.750 0.670 2.330 0.910 ;
        RECT  2.140 1.430 2.260 1.830 ;
        RECT  1.870 2.550 2.110 3.110 ;
        RECT  1.700 3.390 1.940 4.370 ;
        RECT  1.710 2.870 1.870 3.110 ;
        RECT  0.570 3.390 1.700 3.630 ;
        RECT  0.400 1.270 0.570 1.670 ;
        RECT  0.400 2.940 0.570 3.630 ;
        RECT  0.160 1.270 0.400 3.630 ;
    END
END SDFFSXL

MACRO SDFFSX4
    CLASS CORE ;
    FOREIGN SDFFSX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSXL ;
    SIZE 21.780 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.370 4.060 7.990 4.380 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.390 2.020 3.500 2.640 ;
        RECT  3.500 2.020 3.850 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 1.700 1.870 2.260 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.590 1.820 18.860 3.220 ;
        RECT  18.860 1.580 18.870 3.220 ;
        RECT  18.870 1.380 19.030 3.220 ;
        RECT  19.030 1.380 19.270 3.160 ;
        RECT  19.270 1.580 19.280 3.160 ;
        RECT  19.280 2.750 19.330 3.150 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  19.910 1.820 20.200 3.220 ;
        RECT  20.200 1.580 20.210 3.220 ;
        RECT  20.210 1.380 20.470 3.220 ;
        RECT  20.470 1.380 20.610 3.150 ;
        RECT  20.610 1.580 20.620 3.150 ;
        RECT  20.620 2.750 20.870 3.150 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.380 1.760 4.780 2.160 ;
        RECT  4.780 1.830 5.080 2.090 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.690 2.180 0.760 2.640 ;
        RECT  0.760 2.170 1.170 2.660 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.210 5.440 ;
        RECT  0.210 4.480 0.610 5.440 ;
        RECT  0.610 4.640 3.440 5.440 ;
        RECT  3.440 4.110 3.680 5.440 ;
        RECT  3.680 4.640 6.860 5.440 ;
        RECT  6.860 4.170 7.100 5.440 ;
        RECT  7.100 4.640 8.310 5.440 ;
        RECT  8.310 4.260 8.320 5.440 ;
        RECT  8.320 4.060 8.720 5.440 ;
        RECT  8.720 4.260 8.730 5.440 ;
        RECT  8.730 4.640 9.660 5.440 ;
        RECT  9.660 4.270 9.670 5.440 ;
        RECT  9.670 4.070 10.070 5.440 ;
        RECT  10.070 4.270 10.080 5.440 ;
        RECT  10.080 4.640 12.210 5.440 ;
        RECT  12.210 3.830 12.220 5.440 ;
        RECT  12.220 3.630 12.620 5.440 ;
        RECT  12.620 3.830 12.630 5.440 ;
        RECT  12.630 4.640 13.870 5.440 ;
        RECT  13.870 4.080 14.270 5.440 ;
        RECT  14.270 4.640 15.380 5.440 ;
        RECT  15.380 3.490 15.780 5.440 ;
        RECT  15.780 4.640 16.900 5.440 ;
        RECT  16.900 4.480 17.300 5.440 ;
        RECT  17.300 4.640 18.280 5.440 ;
        RECT  18.280 4.210 18.290 5.440 ;
        RECT  18.290 4.010 18.690 5.440 ;
        RECT  18.690 4.210 18.700 5.440 ;
        RECT  18.700 4.640 19.690 5.440 ;
        RECT  19.690 4.210 19.700 5.440 ;
        RECT  19.700 4.010 20.100 5.440 ;
        RECT  20.100 4.210 20.110 5.440 ;
        RECT  20.110 4.640 21.100 5.440 ;
        RECT  21.100 4.210 21.110 5.440 ;
        RECT  21.110 4.010 21.510 5.440 ;
        RECT  21.510 4.210 21.520 5.440 ;
        RECT  21.520 4.640 21.780 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.180 0.400 ;
        RECT  1.180 -0.400 1.580 0.560 ;
        RECT  1.580 -0.400 3.340 0.400 ;
        RECT  3.340 -0.400 3.740 0.560 ;
        RECT  3.740 -0.400 6.890 0.400 ;
        RECT  6.890 -0.400 6.900 1.000 ;
        RECT  6.900 -0.400 7.300 1.120 ;
        RECT  7.300 -0.400 7.310 1.000 ;
        RECT  7.310 -0.400 9.790 0.400 ;
        RECT  9.790 -0.400 9.800 1.160 ;
        RECT  9.800 -0.400 10.200 1.280 ;
        RECT  10.200 -0.400 10.210 1.160 ;
        RECT  10.210 -0.400 12.310 0.400 ;
        RECT  12.310 -0.400 12.710 1.020 ;
        RECT  12.710 -0.400 14.100 0.400 ;
        RECT  14.100 -0.400 14.500 0.560 ;
        RECT  14.500 -0.400 16.620 0.400 ;
        RECT  16.620 -0.400 17.020 0.560 ;
        RECT  17.020 -0.400 18.160 0.400 ;
        RECT  18.160 -0.400 18.170 0.900 ;
        RECT  18.170 -0.400 18.570 1.100 ;
        RECT  18.570 -0.400 18.580 0.900 ;
        RECT  18.580 -0.400 19.530 0.400 ;
        RECT  19.530 -0.400 19.540 0.900 ;
        RECT  19.540 -0.400 19.940 1.100 ;
        RECT  19.940 -0.400 19.950 0.900 ;
        RECT  19.950 -0.400 20.840 0.400 ;
        RECT  20.840 -0.400 20.850 0.900 ;
        RECT  20.850 -0.400 21.250 1.100 ;
        RECT  21.250 -0.400 21.260 0.900 ;
        RECT  21.260 -0.400 21.780 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  21.120 2.070 21.360 3.730 ;
        RECT  18.320 3.490 21.120 3.730 ;
        RECT  18.080 1.390 18.320 3.730 ;
        RECT  17.810 1.390 18.080 1.630 ;
        RECT  17.420 2.750 18.080 3.150 ;
        RECT  17.410 1.200 17.810 1.630 ;
        RECT  17.560 2.050 17.800 2.450 ;
        RECT  16.420 2.050 17.560 2.440 ;
        RECT  16.190 2.050 16.420 3.810 ;
        RECT  16.180 1.550 16.190 3.810 ;
        RECT  15.950 1.550 16.180 2.290 ;
        RECT  14.980 2.860 16.180 3.100 ;
        RECT  15.750 1.550 15.950 1.790 ;
        RECT  15.350 0.890 15.750 1.790 ;
        RECT  15.290 2.220 15.690 2.620 ;
        RECT  14.220 1.550 15.350 1.790 ;
        RECT  13.520 2.380 15.290 2.620 ;
        RECT  14.740 2.860 14.980 3.810 ;
        RECT  13.980 1.550 14.220 2.140 ;
        RECT  13.820 1.900 13.980 2.140 ;
        RECT  13.500 2.380 13.520 3.210 ;
        RECT  13.280 1.500 13.500 3.210 ;
        RECT  13.260 1.500 13.280 2.620 ;
        RECT  11.260 2.970 13.280 3.210 ;
        RECT  12.130 1.500 13.260 1.740 ;
        RECT  12.630 2.170 12.870 2.570 ;
        RECT  11.650 2.250 12.630 2.490 ;
        RECT  11.890 1.240 12.130 1.740 ;
        RECT  11.420 1.240 11.890 1.480 ;
        RECT  11.410 1.720 11.650 2.490 ;
        RECT  10.980 1.110 11.420 1.480 ;
        RECT  10.240 1.800 11.410 2.040 ;
        RECT  11.020 2.970 11.260 3.470 ;
        RECT  10.740 2.380 11.050 2.620 ;
        RECT  10.500 2.380 10.740 3.830 ;
        RECT  9.240 3.590 10.500 3.830 ;
        RECT  10.110 1.520 10.240 2.040 ;
        RECT  9.870 1.520 10.110 3.270 ;
        RECT  9.240 1.520 9.870 1.760 ;
        RECT  9.140 3.030 9.870 3.270 ;
        RECT  9.390 2.240 9.630 2.640 ;
        RECT  8.860 2.320 9.390 2.560 ;
        RECT  9.000 0.670 9.240 1.760 ;
        RECT  9.000 3.550 9.240 4.130 ;
        RECT  8.860 0.670 9.000 1.070 ;
        RECT  6.580 3.550 9.000 3.790 ;
        RECT  8.620 2.000 8.860 3.270 ;
        RECT  8.500 2.000 8.620 2.240 ;
        RECT  7.400 3.030 8.620 3.270 ;
        RECT  8.260 0.930 8.500 2.240 ;
        RECT  7.930 2.480 8.340 2.720 ;
        RECT  7.690 1.400 7.930 2.720 ;
        RECT  6.200 1.400 7.690 1.640 ;
        RECT  7.160 2.090 7.400 3.270 ;
        RECT  7.080 2.090 7.160 2.330 ;
        RECT  6.840 1.930 7.080 2.330 ;
        RECT  6.340 3.550 6.580 4.290 ;
        RECT  5.540 4.050 6.340 4.290 ;
        RECT  6.060 1.360 6.200 3.130 ;
        RECT  5.960 1.360 6.060 3.760 ;
        RECT  5.560 0.990 5.960 1.640 ;
        RECT  5.820 2.890 5.960 3.760 ;
        RECT  5.540 1.990 5.680 2.610 ;
        RECT  5.440 1.990 5.540 4.290 ;
        RECT  5.300 2.370 5.440 4.290 ;
        RECT  4.440 4.050 5.300 4.290 ;
        RECT  5.000 0.890 5.080 1.290 ;
        RECT  4.780 3.070 5.020 3.620 ;
        RECT  4.680 0.860 5.000 1.290 ;
        RECT  2.640 3.070 4.780 3.310 ;
        RECT  2.380 0.860 4.680 1.100 ;
        RECT  4.200 3.590 4.440 4.290 ;
        RECT  3.160 3.590 4.200 3.830 ;
        RECT  2.380 1.380 4.040 1.620 ;
        RECT  2.920 3.590 3.160 4.370 ;
        RECT  2.380 2.540 2.930 2.780 ;
        RECT  1.690 4.130 2.920 4.370 ;
        RECT  2.400 3.070 2.640 3.850 ;
        RECT  2.230 3.610 2.400 3.850 ;
        RECT  1.980 0.670 2.380 1.100 ;
        RECT  2.140 1.380 2.380 2.780 ;
        RECT  2.070 2.540 2.140 2.780 ;
        RECT  1.830 2.540 2.070 3.110 ;
        RECT  1.650 2.870 1.830 3.110 ;
        RECT  1.450 3.390 1.690 4.370 ;
        RECT  0.570 3.390 1.450 3.630 ;
        RECT  0.410 1.240 0.570 1.640 ;
        RECT  0.410 2.930 0.570 3.630 ;
        RECT  0.330 1.240 0.410 3.630 ;
        RECT  0.170 1.240 0.330 3.330 ;
    END
END SDFFSX4

MACRO SDFFSX2
    CLASS CORE ;
    FOREIGN SDFFSX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.800 1.830 6.910 2.090 ;
        RECT  6.910 1.830 7.060 2.100 ;
        RECT  7.060 1.840 7.150 2.100 ;
        RECT  7.150 1.860 7.350 2.100 ;
        RECT  7.350 1.860 7.590 2.400 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.160 2.010 3.560 2.650 ;
        RECT  3.560 2.390 3.760 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.740 1.950 2.180 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.150 2.790 15.180 3.190 ;
        RECT  15.180 2.600 15.190 3.190 ;
        RECT  15.030 0.670 15.190 0.910 ;
        RECT  15.190 0.670 15.430 3.190 ;
        RECT  15.430 2.390 15.630 3.190 ;
        RECT  15.630 2.390 15.640 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.040 1.270 16.150 1.530 ;
        RECT  16.150 1.260 16.590 1.540 ;
        RECT  16.590 0.700 16.610 1.680 ;
        RECT  16.590 3.130 16.670 4.110 ;
        RECT  16.610 0.700 16.670 1.820 ;
        RECT  16.670 0.700 16.910 4.110 ;
        RECT  16.910 3.130 16.990 4.110 ;
        RECT  16.910 0.700 16.990 1.840 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.530 1.380 4.730 1.620 ;
        RECT  4.730 1.260 5.170 1.630 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.730 2.120 1.170 2.660 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.480 5.440 ;
        RECT  0.480 4.480 0.880 5.440 ;
        RECT  0.880 4.640 3.400 5.440 ;
        RECT  3.400 4.110 3.640 5.440 ;
        RECT  3.640 4.640 6.830 5.440 ;
        RECT  6.830 4.480 7.230 5.440 ;
        RECT  7.230 4.640 8.350 5.440 ;
        RECT  8.350 4.240 8.360 5.440 ;
        RECT  8.360 4.120 8.760 5.440 ;
        RECT  8.760 4.240 8.770 5.440 ;
        RECT  8.770 4.640 9.750 5.440 ;
        RECT  9.750 4.220 9.760 5.440 ;
        RECT  9.760 4.020 10.160 5.440 ;
        RECT  10.160 4.220 10.170 5.440 ;
        RECT  10.170 4.640 12.140 5.440 ;
        RECT  12.140 3.780 12.150 5.440 ;
        RECT  12.150 3.580 12.550 5.440 ;
        RECT  12.550 3.780 12.560 5.440 ;
        RECT  12.560 4.640 13.720 5.440 ;
        RECT  13.720 4.480 14.120 5.440 ;
        RECT  14.120 4.640 15.820 5.440 ;
        RECT  15.820 4.290 15.830 5.440 ;
        RECT  15.830 4.090 16.230 5.440 ;
        RECT  16.230 4.290 16.240 5.440 ;
        RECT  16.240 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.180 0.400 ;
        RECT  1.180 -0.400 1.580 0.560 ;
        RECT  1.580 -0.400 3.450 0.400 ;
        RECT  3.450 -0.400 3.850 0.560 ;
        RECT  3.850 -0.400 7.060 0.400 ;
        RECT  7.060 -0.400 7.070 0.910 ;
        RECT  7.070 -0.400 7.470 1.030 ;
        RECT  7.470 -0.400 7.480 0.910 ;
        RECT  7.480 -0.400 9.550 0.400 ;
        RECT  9.550 -0.400 9.790 1.110 ;
        RECT  9.790 -0.400 12.090 0.400 ;
        RECT  12.090 -0.400 12.490 0.560 ;
        RECT  12.490 -0.400 13.880 0.400 ;
        RECT  13.880 -0.400 14.280 0.560 ;
        RECT  14.280 -0.400 15.820 0.400 ;
        RECT  15.820 -0.400 15.830 0.720 ;
        RECT  15.830 -0.400 16.230 0.920 ;
        RECT  16.230 -0.400 16.240 0.720 ;
        RECT  16.240 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.310 2.220 16.390 2.620 ;
        RECT  16.070 2.220 16.310 3.710 ;
        RECT  14.870 3.470 16.070 3.710 ;
        RECT  14.870 1.330 14.910 1.730 ;
        RECT  14.630 1.330 14.870 3.710 ;
        RECT  14.510 1.330 14.630 1.730 ;
        RECT  14.330 3.120 14.630 3.710 ;
        RECT  13.590 2.020 14.350 2.420 ;
        RECT  13.350 1.160 13.590 3.150 ;
        RECT  13.010 1.160 13.350 1.400 ;
        RECT  13.310 2.910 13.350 3.150 ;
        RECT  12.910 2.910 13.310 3.380 ;
        RECT  12.670 1.890 13.070 2.400 ;
        RECT  12.610 1.000 13.010 1.400 ;
        RECT  12.350 2.910 12.910 3.150 ;
        RECT  11.670 1.890 12.670 2.130 ;
        RECT  12.190 1.160 12.610 1.400 ;
        RECT  12.110 2.410 12.350 3.150 ;
        RECT  11.790 1.160 12.190 1.610 ;
        RECT  11.950 2.410 12.110 2.650 ;
        RECT  11.510 1.890 11.670 3.940 ;
        RECT  11.430 1.300 11.510 3.940 ;
        RECT  11.270 1.300 11.430 2.130 ;
        RECT  11.070 1.300 11.270 1.540 ;
        RECT  10.860 3.500 11.100 4.290 ;
        RECT  10.830 1.140 11.070 1.540 ;
        RECT  10.550 1.820 10.930 2.060 ;
        RECT  9.480 3.500 10.860 3.740 ;
        RECT  10.310 1.390 10.550 3.120 ;
        RECT  9.260 1.390 10.310 1.630 ;
        RECT  9.240 2.880 10.310 3.120 ;
        RECT  9.790 2.150 10.030 2.550 ;
        RECT  8.960 2.230 9.790 2.470 ;
        RECT  9.240 3.500 9.480 3.840 ;
        RECT  9.020 0.670 9.260 1.630 ;
        RECT  6.540 3.600 9.240 3.840 ;
        RECT  8.020 0.670 9.020 0.910 ;
        RECT  8.730 1.990 8.960 3.310 ;
        RECT  8.720 1.430 8.730 3.310 ;
        RECT  8.490 1.430 8.720 2.230 ;
        RECT  6.730 3.070 8.720 3.310 ;
        RECT  8.070 2.510 8.440 2.750 ;
        RECT  7.830 1.310 8.070 2.750 ;
        RECT  6.210 1.310 7.830 1.550 ;
        RECT  6.490 2.430 6.730 3.310 ;
        RECT  6.300 3.600 6.540 4.250 ;
        RECT  5.500 4.010 6.300 4.250 ;
        RECT  6.020 0.850 6.210 3.320 ;
        RECT  5.970 0.850 6.020 3.580 ;
        RECT  5.670 0.850 5.970 1.250 ;
        RECT  5.780 3.080 5.970 3.580 ;
        RECT  5.260 2.020 5.500 4.250 ;
        RECT  3.120 3.590 5.260 3.830 ;
        RECT  4.370 0.750 5.190 0.990 ;
        RECT  4.740 2.910 4.980 3.310 ;
        RECT  2.600 3.070 4.740 3.310 ;
        RECT  4.130 0.750 4.370 1.100 ;
        RECT  2.460 1.380 4.170 1.620 ;
        RECT  2.510 0.860 4.130 1.100 ;
        RECT  2.880 3.590 3.120 4.370 ;
        RECT  1.880 4.130 2.880 4.370 ;
        RECT  2.460 2.470 2.820 2.710 ;
        RECT  2.360 3.070 2.600 3.850 ;
        RECT  2.110 0.670 2.510 1.100 ;
        RECT  2.220 1.380 2.460 2.710 ;
        RECT  2.120 3.610 2.360 3.850 ;
        RECT  2.080 2.470 2.220 2.710 ;
        RECT  1.840 2.470 2.080 3.190 ;
        RECT  1.640 3.540 1.880 4.370 ;
        RECT  1.680 2.790 1.840 3.190 ;
        RECT  0.600 3.540 1.640 3.780 ;
        RECT  0.520 1.270 0.920 1.670 ;
        RECT  0.460 2.930 0.600 3.780 ;
        RECT  0.460 1.430 0.520 1.670 ;
        RECT  0.360 1.430 0.460 3.780 ;
        RECT  0.220 1.430 0.360 3.330 ;
        RECT  0.200 2.930 0.220 3.330 ;
    END
END SDFFSX2

MACRO SDFFSX1
    CLASS CORE ;
    FOREIGN SDFFSX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFSXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  12.740 4.070 12.750 4.330 ;
        RECT  12.750 3.900 13.000 4.330 ;
        RECT  13.000 3.900 13.080 4.140 ;
        RECT  13.080 3.740 13.320 4.140 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.350 2.160 3.410 2.640 ;
        RECT  3.410 2.150 3.810 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.330 1.820 1.870 2.170 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.290 0.670 14.690 1.100 ;
        RECT  14.340 3.650 14.720 4.050 ;
        RECT  14.720 3.510 14.970 4.050 ;
        RECT  14.970 3.510 14.980 3.770 ;
        RECT  14.980 3.520 15.410 3.760 ;
        RECT  14.690 0.860 15.410 1.100 ;
        RECT  15.410 0.860 15.650 3.760 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.930 1.320 15.950 1.720 ;
        RECT  15.950 1.320 16.040 1.820 ;
        RECT  15.930 2.980 16.050 3.380 ;
        RECT  16.040 1.320 16.050 2.090 ;
        RECT  16.050 1.320 16.290 3.380 ;
        RECT  16.290 1.320 16.300 2.090 ;
        RECT  16.290 2.980 16.330 3.380 ;
        RECT  16.300 1.320 16.330 1.960 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.110 1.440 4.160 1.840 ;
        RECT  4.160 1.440 4.420 2.090 ;
        RECT  4.420 1.440 4.510 1.840 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.700 2.180 0.780 2.580 ;
        RECT  0.780 2.180 0.790 3.200 ;
        RECT  0.790 2.170 0.860 3.200 ;
        RECT  0.860 2.170 1.050 3.210 ;
        RECT  1.050 2.950 1.120 3.210 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.200 5.440 ;
        RECT  0.200 4.480 0.600 5.440 ;
        RECT  0.600 4.640 3.430 5.440 ;
        RECT  3.430 4.070 3.670 5.440 ;
        RECT  3.670 4.640 6.860 5.440 ;
        RECT  6.860 4.480 7.260 5.440 ;
        RECT  7.260 4.640 8.380 5.440 ;
        RECT  8.380 4.290 8.390 5.440 ;
        RECT  8.390 4.090 8.790 5.440 ;
        RECT  8.790 4.290 8.800 5.440 ;
        RECT  8.800 4.640 9.530 5.440 ;
        RECT  9.530 4.290 9.540 5.440 ;
        RECT  9.540 4.090 9.940 5.440 ;
        RECT  9.940 4.290 9.950 5.440 ;
        RECT  9.950 4.640 11.930 5.440 ;
        RECT  11.930 3.790 11.940 5.440 ;
        RECT  11.940 3.590 12.340 5.440 ;
        RECT  12.340 3.790 12.350 5.440 ;
        RECT  12.350 4.640 13.590 5.440 ;
        RECT  13.520 3.060 13.590 3.460 ;
        RECT  13.590 3.050 14.010 5.440 ;
        RECT  14.010 4.640 15.130 5.440 ;
        RECT  15.130 4.480 15.530 5.440 ;
        RECT  15.530 4.640 16.500 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 2.920 0.400 ;
        RECT  2.920 -0.400 3.320 0.560 ;
        RECT  3.320 -0.400 6.470 0.400 ;
        RECT  6.470 -0.400 6.480 0.880 ;
        RECT  6.480 -0.400 6.880 1.000 ;
        RECT  6.880 -0.400 6.890 0.880 ;
        RECT  6.890 -0.400 9.130 0.400 ;
        RECT  9.130 -0.400 9.370 0.950 ;
        RECT  9.370 -0.400 11.630 0.400 ;
        RECT  11.630 -0.400 12.030 0.560 ;
        RECT  12.030 -0.400 13.520 0.400 ;
        RECT  13.520 -0.400 13.530 0.670 ;
        RECT  13.530 -0.400 13.930 0.870 ;
        RECT  13.930 -0.400 13.940 0.670 ;
        RECT  13.940 -0.400 15.100 0.400 ;
        RECT  15.100 -0.400 15.500 0.560 ;
        RECT  15.500 -0.400 16.500 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.800 2.080 15.130 2.480 ;
        RECT  14.560 1.380 14.800 3.230 ;
        RECT  14.350 1.380 14.560 1.780 ;
        RECT  14.400 2.990 14.560 3.230 ;
        RECT  13.820 2.110 14.220 2.510 ;
        RECT  13.160 2.190 13.820 2.430 ;
        RECT  12.920 1.630 13.160 3.430 ;
        RECT  12.650 1.630 12.920 1.870 ;
        RECT  12.760 3.030 12.920 3.430 ;
        RECT  12.250 1.160 12.650 1.870 ;
        RECT  12.380 2.350 12.620 2.750 ;
        RECT  11.280 2.430 12.380 2.670 ;
        RECT  12.000 1.630 12.250 1.870 ;
        RECT  11.600 1.630 12.000 2.030 ;
        RECT  11.040 1.230 11.280 3.920 ;
        RECT  10.390 1.230 11.040 1.470 ;
        RECT  10.900 3.520 11.040 3.920 ;
        RECT  10.380 2.520 10.620 3.810 ;
        RECT  10.100 1.840 10.480 2.080 ;
        RECT  6.570 3.570 10.380 3.810 ;
        RECT  9.860 1.230 10.100 2.920 ;
        RECT  8.810 1.230 9.860 1.470 ;
        RECT  9.590 2.680 9.860 2.920 ;
        RECT  9.350 2.680 9.590 3.180 ;
        RECT  9.340 1.750 9.580 2.150 ;
        RECT  9.050 1.830 9.340 2.070 ;
        RECT  8.810 1.830 9.050 3.290 ;
        RECT  8.570 0.670 8.810 1.470 ;
        RECT  8.290 1.830 8.810 2.070 ;
        RECT  7.110 3.050 8.810 3.290 ;
        RECT  7.160 0.670 8.570 0.910 ;
        RECT  8.050 1.370 8.290 2.070 ;
        RECT  7.950 2.350 8.190 2.770 ;
        RECT  7.630 2.350 7.950 2.590 ;
        RECT  7.390 1.280 7.630 2.590 ;
        RECT  6.050 1.280 7.390 1.520 ;
        RECT  6.870 2.130 7.110 3.290 ;
        RECT  6.810 2.130 6.870 2.370 ;
        RECT  6.570 1.970 6.810 2.370 ;
        RECT  6.330 3.570 6.570 4.090 ;
        RECT  5.530 3.850 6.330 4.090 ;
        RECT  5.810 1.010 6.050 3.560 ;
        RECT  5.540 1.010 5.810 1.250 ;
        RECT  5.140 0.850 5.540 1.250 ;
        RECT  5.290 1.690 5.530 4.090 ;
        RECT  5.160 1.690 5.290 1.930 ;
        RECT  4.480 3.850 5.290 4.090 ;
        RECT  4.920 1.530 5.160 1.930 ;
        RECT  4.770 3.030 5.010 3.500 ;
        RECT  2.570 3.030 4.770 3.270 ;
        RECT  4.260 0.750 4.660 1.150 ;
        RECT  4.240 3.550 4.480 4.090 ;
        RECT  1.980 0.860 4.260 1.100 ;
        RECT  3.090 3.550 4.240 3.790 ;
        RECT  2.380 1.380 3.620 1.620 ;
        RECT  2.850 3.550 3.090 4.370 ;
        RECT  1.690 4.130 2.850 4.370 ;
        RECT  2.330 3.030 2.570 3.850 ;
        RECT  2.140 1.380 2.380 2.680 ;
        RECT  2.170 3.610 2.330 3.850 ;
        RECT  2.050 2.440 2.140 2.680 ;
        RECT  1.810 2.440 2.050 3.190 ;
        RECT  1.570 0.670 1.980 1.100 ;
        RECT  1.650 2.790 1.810 3.190 ;
        RECT  1.450 3.650 1.690 4.370 ;
        RECT  0.490 3.650 1.450 3.890 ;
        RECT  0.400 1.270 0.570 1.670 ;
        RECT  0.400 2.860 0.490 3.890 ;
        RECT  0.250 1.270 0.400 3.890 ;
        RECT  0.160 1.270 0.250 3.280 ;
    END
END SDFFSX1

MACRO SDFFRHQXL
    CLASS CORE ;
    FOREIGN SDFFRHQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.110 2.020 3.500 2.640 ;
        RECT  3.500 2.020 3.510 2.650 ;
        RECT  3.510 2.390 3.760 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.470 1.830 1.870 2.280 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  14.490 2.910 15.070 3.260 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.350 1.000 15.590 1.400 ;
        RECT  15.920 3.600 15.990 4.000 ;
        RECT  15.990 2.950 16.090 4.010 ;
        RECT  15.590 1.160 16.090 1.400 ;
        RECT  16.090 1.160 16.330 4.010 ;
        RECT  16.330 2.950 16.340 4.010 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.110 1.830 4.510 2.350 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.100 0.780 2.500 ;
        RECT  0.780 2.100 0.860 2.640 ;
        RECT  0.860 2.080 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.750 5.440 ;
        RECT  0.750 3.770 0.990 5.440 ;
        RECT  0.990 4.640 3.370 5.440 ;
        RECT  3.370 4.110 3.610 5.440 ;
        RECT  3.610 4.640 6.460 5.440 ;
        RECT  6.460 4.080 7.440 5.440 ;
        RECT  7.440 4.640 9.410 5.440 ;
        RECT  9.410 4.480 9.810 5.440 ;
        RECT  9.810 4.640 12.560 5.440 ;
        RECT  12.560 4.480 12.960 5.440 ;
        RECT  13.770 3.310 14.170 3.770 ;
        RECT  12.960 4.640 14.700 5.440 ;
        RECT  14.170 3.530 14.700 3.770 ;
        RECT  14.700 3.530 14.940 5.440 ;
        RECT  14.940 3.780 15.100 5.440 ;
        RECT  15.100 4.640 16.500 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.050 0.400 ;
        RECT  1.050 -0.400 1.450 0.560 ;
        RECT  1.450 -0.400 3.130 0.400 ;
        RECT  3.130 -0.400 3.530 0.560 ;
        RECT  3.530 -0.400 6.550 0.400 ;
        RECT  6.550 -0.400 6.950 1.440 ;
        RECT  6.950 1.200 8.090 1.440 ;
        RECT  8.090 1.200 8.490 1.830 ;
        RECT  6.950 -0.400 9.300 0.400 ;
        RECT  9.300 -0.400 9.540 1.160 ;
        RECT  9.540 -0.400 12.200 0.400 ;
        RECT  12.200 -0.400 12.600 0.560 ;
        RECT  12.600 -0.400 13.820 0.400 ;
        RECT  13.820 -0.400 14.800 0.560 ;
        RECT  14.800 -0.400 15.940 0.400 ;
        RECT  15.940 -0.400 16.340 0.560 ;
        RECT  16.340 -0.400 16.500 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  15.570 1.680 15.810 2.080 ;
        RECT  15.340 2.360 15.580 2.810 ;
        RECT  15.070 1.680 15.570 1.920 ;
        RECT  14.370 2.360 15.340 2.600 ;
        RECT  14.830 0.910 15.070 1.920 ;
        RECT  12.210 0.910 14.830 1.150 ;
        RECT  13.970 1.600 14.370 2.600 ;
        RECT  13.490 4.130 14.220 4.370 ;
        RECT  13.930 2.360 13.970 2.600 ;
        RECT  13.530 2.360 13.930 2.760 ;
        RECT  13.490 2.520 13.530 2.760 ;
        RECT  13.250 2.520 13.490 4.370 ;
        RECT  12.790 1.480 13.310 1.720 ;
        RECT  8.450 3.940 13.250 4.180 ;
        RECT  12.790 3.210 12.950 3.610 ;
        RECT  12.550 1.480 12.790 3.610 ;
        RECT  12.430 2.630 12.550 3.610 ;
        RECT  12.150 0.910 12.210 2.350 ;
        RECT  11.970 0.910 12.150 3.660 ;
        RECT  11.180 0.910 11.970 1.150 ;
        RECT  11.910 2.110 11.970 3.660 ;
        RECT  11.230 3.420 11.910 3.660 ;
        RECT  11.330 1.660 11.560 1.900 ;
        RECT  11.090 1.660 11.330 3.140 ;
        RECT  10.940 0.910 11.180 1.350 ;
        RECT  10.810 3.410 10.870 3.650 ;
        RECT  10.660 1.780 10.810 3.650 ;
        RECT  10.570 1.060 10.660 3.650 ;
        RECT  10.420 1.060 10.570 2.020 ;
        RECT  10.470 3.410 10.570 3.650 ;
        RECT  10.100 1.060 10.420 1.300 ;
        RECT  10.140 2.300 10.290 2.700 ;
        RECT  9.900 1.580 10.140 3.660 ;
        RECT  9.020 1.580 9.900 1.820 ;
        RECT  9.070 3.420 9.900 3.660 ;
        RECT  9.330 2.170 9.570 2.600 ;
        RECT  7.770 2.170 9.330 2.410 ;
        RECT  8.780 0.680 9.020 1.820 ;
        RECT  7.230 0.680 8.780 0.920 ;
        RECT  8.210 2.690 8.450 4.180 ;
        RECT  8.050 2.690 8.210 2.930 ;
        RECT  7.610 2.030 7.770 3.550 ;
        RECT  7.530 1.720 7.610 3.550 ;
        RECT  7.210 1.720 7.530 2.270 ;
        RECT  7.410 3.310 7.530 3.550 ;
        RECT  7.170 3.310 7.410 3.710 ;
        RECT  6.990 2.550 7.230 2.950 ;
        RECT  6.510 2.030 7.210 2.270 ;
        RECT  5.930 2.710 6.990 2.950 ;
        RECT  6.270 2.000 6.510 2.400 ;
        RECT  5.690 0.670 5.930 2.950 ;
        RECT  5.030 3.940 5.930 4.180 ;
        RECT  5.210 0.670 5.690 0.910 ;
        RECT  5.550 2.710 5.690 2.950 ;
        RECT  5.310 2.710 5.550 3.560 ;
        RECT  5.030 1.940 5.350 2.340 ;
        RECT  4.790 1.940 5.030 4.180 ;
        RECT  4.470 0.740 4.870 1.140 ;
        RECT  2.550 3.070 4.790 3.310 ;
        RECT  4.270 3.590 4.510 4.360 ;
        RECT  2.190 0.860 4.470 1.100 ;
        RECT  3.070 3.590 4.270 3.830 ;
        RECT  2.380 1.380 3.740 1.620 ;
        RECT  2.830 3.590 3.070 4.230 ;
        RECT  2.170 3.990 2.830 4.230 ;
        RECT  2.380 2.550 2.680 2.790 ;
        RECT  2.310 3.070 2.550 3.710 ;
        RECT  2.140 1.380 2.380 2.790 ;
        RECT  1.510 3.470 2.310 3.710 ;
        RECT  1.790 0.670 2.190 1.100 ;
        RECT  2.030 2.550 2.140 2.790 ;
        RECT  1.790 2.550 2.030 3.190 ;
        RECT  1.270 2.950 1.510 3.710 ;
        RECT  0.490 2.950 1.270 3.190 ;
        RECT  0.400 1.260 0.490 1.660 ;
        RECT  0.400 2.790 0.490 3.190 ;
        RECT  0.160 1.260 0.400 3.190 ;
    END
END SDFFRHQXL

MACRO SDFFRHQX4
    CLASS CORE ;
    FOREIGN SDFFRHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFRHQXL ;
    SIZE 24.420 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.760 2.940 3.310 3.340 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.780 1.960 2.940 2.520 ;
        RECT  2.940 1.960 3.180 2.610 ;
        RECT  3.180 2.370 3.500 2.610 ;
        RECT  3.500 2.370 3.760 2.650 ;
        RECT  3.760 2.370 4.320 2.610 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  17.800 1.630 18.280 2.120 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.340 0.730 21.740 1.710 ;
        RECT  21.390 2.960 21.790 3.940 ;
        RECT  21.790 2.960 22.110 3.220 ;
        RECT  22.110 2.980 22.770 3.220 ;
        RECT  21.740 1.460 22.860 1.700 ;
        RECT  22.770 2.940 23.210 3.220 ;
        RECT  22.860 0.730 23.210 1.710 ;
        RECT  23.210 0.730 23.260 3.220 ;
        RECT  23.260 1.450 23.650 3.220 ;
        RECT  23.650 2.940 23.830 3.220 ;
        RECT  23.830 2.940 24.100 3.930 ;
        RECT  24.100 2.950 24.230 3.930 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 2.950 4.370 3.210 ;
        RECT  4.370 2.950 4.420 3.330 ;
        RECT  4.420 2.960 4.770 3.330 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 1.970 0.860 2.640 ;
        RECT  0.860 1.970 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.980 5.440 ;
        RECT  0.980 4.480 1.380 5.440 ;
        RECT  1.380 4.640 6.800 5.440 ;
        RECT  6.800 4.480 7.200 5.440 ;
        RECT  7.200 4.640 8.590 5.440 ;
        RECT  8.590 4.480 8.990 5.440 ;
        RECT  8.990 4.640 10.240 5.440 ;
        RECT  10.240 4.010 10.480 5.440 ;
        RECT  10.480 4.640 11.780 5.440 ;
        RECT  11.780 4.480 12.180 5.440 ;
        RECT  12.180 4.640 17.070 5.440 ;
        RECT  17.070 4.190 17.310 5.440 ;
        RECT  17.310 4.640 18.640 5.440 ;
        RECT  18.640 4.480 19.040 5.440 ;
        RECT  19.040 4.640 20.250 5.440 ;
        RECT  20.250 3.080 20.490 5.440 ;
        RECT  20.490 4.640 22.600 5.440 ;
        RECT  22.600 3.930 22.610 5.440 ;
        RECT  22.610 3.730 23.010 5.440 ;
        RECT  23.010 3.930 23.020 5.440 ;
        RECT  23.020 4.640 24.420 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        RECT  0.990 -0.400 1.390 0.560 ;
        RECT  1.390 -0.400 3.810 0.400 ;
        RECT  3.810 -0.400 4.210 0.560 ;
        RECT  4.210 -0.400 6.960 0.400 ;
        RECT  6.960 -0.400 6.970 0.800 ;
        RECT  6.970 -0.400 7.370 1.000 ;
        RECT  7.370 -0.400 7.380 0.800 ;
        RECT  7.380 -0.400 8.450 0.400 ;
        RECT  8.450 -0.400 8.630 1.470 ;
        RECT  8.630 -0.400 8.690 1.630 ;
        RECT  8.690 1.230 8.870 1.630 ;
        RECT  8.690 -0.400 10.050 0.400 ;
        RECT  10.050 -0.400 10.060 1.250 ;
        RECT  10.060 -0.400 10.460 1.450 ;
        RECT  10.460 -0.400 10.470 1.250 ;
        RECT  10.470 -0.400 11.570 0.400 ;
        RECT  11.570 -0.400 11.580 1.150 ;
        RECT  11.580 -0.400 11.980 1.270 ;
        RECT  11.980 -0.400 11.990 1.150 ;
        RECT  11.990 -0.400 17.290 0.400 ;
        RECT  17.290 -0.400 17.300 1.020 ;
        RECT  17.300 -0.400 17.700 1.220 ;
        RECT  17.700 -0.400 17.710 1.020 ;
        RECT  17.710 -0.400 18.880 0.400 ;
        RECT  18.880 -0.400 19.280 0.560 ;
        RECT  19.280 -0.400 20.660 0.400 ;
        RECT  20.660 -0.400 20.900 1.650 ;
        RECT  20.900 -0.400 22.090 0.400 ;
        RECT  22.090 -0.400 22.100 0.880 ;
        RECT  22.100 -0.400 22.500 1.080 ;
        RECT  22.500 -0.400 22.510 0.880 ;
        RECT  22.510 -0.400 23.610 0.400 ;
        RECT  23.610 -0.400 23.620 0.880 ;
        RECT  23.620 -0.400 24.020 1.080 ;
        RECT  24.020 -0.400 24.030 0.880 ;
        RECT  24.030 -0.400 24.420 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  20.380 2.120 22.770 2.360 ;
        RECT  20.140 0.860 20.380 2.500 ;
        RECT  18.380 0.860 20.140 1.100 ;
        RECT  19.970 2.260 20.140 2.500 ;
        RECT  19.730 2.260 19.970 4.180 ;
        RECT  19.620 1.380 19.860 1.780 ;
        RECT  18.210 3.940 19.730 4.180 ;
        RECT  18.900 1.540 19.620 1.780 ;
        RECT  19.210 2.170 19.450 3.660 ;
        RECT  18.350 3.420 19.210 3.660 ;
        RECT  18.660 1.540 18.900 3.140 ;
        RECT  18.630 2.560 18.660 3.140 ;
        RECT  17.310 2.560 18.630 2.800 ;
        RECT  18.140 0.860 18.380 1.360 ;
        RECT  18.110 3.150 18.350 3.660 ;
        RECT  17.830 3.940 18.210 4.230 ;
        RECT  16.790 3.150 18.110 3.390 ;
        RECT  17.810 3.670 17.830 4.230 ;
        RECT  17.590 3.670 17.810 4.180 ;
        RECT  16.790 3.670 17.590 3.910 ;
        RECT  17.070 2.210 17.310 2.800 ;
        RECT  16.670 2.210 17.070 2.450 ;
        RECT  16.550 2.730 16.790 3.390 ;
        RECT  16.550 3.670 16.790 4.370 ;
        RECT  16.200 2.730 16.550 2.970 ;
        RECT  12.700 4.130 16.550 4.370 ;
        RECT  16.200 1.070 16.360 1.470 ;
        RECT  16.030 3.250 16.270 3.850 ;
        RECT  15.960 0.670 16.200 2.970 ;
        RECT  13.220 3.610 16.030 3.850 ;
        RECT  14.850 0.670 15.960 0.910 ;
        RECT  15.670 2.570 15.960 2.970 ;
        RECT  14.030 2.570 15.670 2.810 ;
        RECT  15.440 1.190 15.600 1.430 ;
        RECT  15.200 1.190 15.440 1.930 ;
        RECT  13.750 3.090 15.250 3.330 ;
        RECT  14.090 1.690 15.200 1.930 ;
        RECT  14.840 0.670 14.850 1.210 ;
        RECT  14.440 0.670 14.840 1.410 ;
        RECT  14.430 0.670 14.440 1.210 ;
        RECT  12.860 0.670 14.430 0.910 ;
        RECT  14.080 1.310 14.090 1.930 ;
        RECT  13.750 1.190 14.080 1.930 ;
        RECT  13.510 1.190 13.750 3.330 ;
        RECT  13.500 1.190 13.510 1.730 ;
        RECT  12.040 2.900 13.510 3.140 ;
        RECT  12.660 1.190 13.500 1.430 ;
        RECT  12.990 1.740 13.230 2.440 ;
        RECT  12.980 3.420 13.220 3.850 ;
        RECT  11.520 2.200 12.990 2.440 ;
        RECT  11.520 3.420 12.980 3.660 ;
        RECT  12.460 3.940 12.700 4.370 ;
        RECT  12.420 1.190 12.660 1.790 ;
        RECT  11.000 3.940 12.460 4.180 ;
        RECT  11.220 1.550 12.420 1.790 ;
        RECT  11.800 2.740 12.040 3.140 ;
        RECT  11.280 2.200 11.520 3.660 ;
        RECT  10.220 2.200 11.280 2.440 ;
        RECT  10.980 1.110 11.220 1.790 ;
        RECT  10.760 3.390 11.000 4.180 ;
        RECT  10.820 1.110 10.980 1.510 ;
        RECT  9.700 3.390 10.760 3.630 ;
        RECT  9.980 1.770 10.220 3.110 ;
        RECT  9.700 1.770 9.980 2.010 ;
        RECT  9.670 3.910 9.910 4.310 ;
        RECT  9.540 1.230 9.700 2.010 ;
        RECT  9.460 2.290 9.700 3.630 ;
        RECT  6.380 3.940 9.670 4.180 ;
        RECT  9.380 0.670 9.540 2.010 ;
        RECT  8.620 2.290 9.460 2.530 ;
        RECT  9.300 0.670 9.380 1.630 ;
        RECT  8.970 0.670 9.300 0.910 ;
        RECT  8.340 2.930 9.180 3.330 ;
        RECT  8.170 1.750 8.340 3.330 ;
        RECT  8.100 1.230 8.170 3.330 ;
        RECT  7.930 1.230 8.100 1.990 ;
        RECT  7.710 3.090 8.100 3.330 ;
        RECT  7.870 1.230 7.930 1.630 ;
        RECT  7.650 2.270 7.820 2.670 ;
        RECT  7.310 3.090 7.710 3.510 ;
        RECT  7.410 2.010 7.650 2.670 ;
        RECT  6.170 2.010 7.410 2.250 ;
        RECT  7.100 3.090 7.310 3.330 ;
        RECT  6.860 2.540 7.100 3.330 ;
        RECT  6.140 2.800 6.380 4.180 ;
        RECT  5.930 0.870 6.170 2.370 ;
        RECT  5.290 3.610 6.140 3.850 ;
        RECT  5.810 2.130 5.930 2.370 ;
        RECT  5.570 2.130 5.810 3.330 ;
        RECT  5.370 1.440 5.610 1.840 ;
        RECT  5.090 0.870 5.490 1.160 ;
        RECT  5.290 1.600 5.370 1.840 ;
        RECT  5.050 1.600 5.290 3.850 ;
        RECT  2.870 0.870 5.090 1.110 ;
        RECT  2.470 3.610 5.050 3.850 ;
        RECT  1.950 4.130 5.030 4.370 ;
        RECT  3.990 1.440 4.390 1.840 ;
        RECT  2.130 1.440 3.990 1.680 ;
        RECT  2.470 0.870 2.870 1.160 ;
        RECT  2.230 3.150 2.470 3.850 ;
        RECT  0.490 3.150 2.230 3.390 ;
        RECT  2.110 1.050 2.130 1.680 ;
        RECT  1.870 1.050 2.110 2.870 ;
        RECT  1.710 3.670 1.950 4.370 ;
        RECT  1.730 1.050 1.870 1.290 ;
        RECT  1.650 2.630 1.870 2.870 ;
        RECT  0.400 1.190 0.570 1.590 ;
        RECT  0.400 3.040 0.490 4.020 ;
        RECT  0.250 1.190 0.400 4.020 ;
        RECT  0.160 1.190 0.250 3.290 ;
    END
END SDFFRHQX4

MACRO SDFFRHQX2
    CLASS CORE ;
    FOREIGN SDFFRHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFRHQXL ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.190 2.020 3.430 2.630 ;
        RECT  3.430 2.390 3.500 2.630 ;
        RECT  3.500 2.390 3.760 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.470 1.830 1.870 2.280 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  16.040 2.950 16.200 3.210 ;
        RECT  16.200 2.740 16.600 3.210 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.570 0.990 17.970 1.390 ;
        RECT  18.010 3.070 18.020 4.050 ;
        RECT  18.020 2.950 18.170 4.050 ;
        RECT  18.170 2.940 18.410 4.050 ;
        RECT  18.410 2.940 18.450 3.180 ;
        RECT  17.970 1.150 18.450 1.390 ;
        RECT  18.450 1.150 18.690 3.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.880 1.740 4.510 2.100 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.180 0.860 2.640 ;
        RECT  0.860 2.180 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.980 5.440 ;
        RECT  0.980 4.190 0.990 5.440 ;
        RECT  0.990 3.990 1.390 5.440 ;
        RECT  1.390 4.190 1.400 5.440 ;
        RECT  1.400 4.640 3.290 5.440 ;
        RECT  3.290 4.110 3.530 5.440 ;
        RECT  3.530 4.640 6.300 5.440 ;
        RECT  6.300 4.160 6.310 5.440 ;
        RECT  6.310 3.960 6.710 5.440 ;
        RECT  6.710 4.160 6.720 5.440 ;
        RECT  6.720 4.640 10.220 5.440 ;
        RECT  10.220 4.480 10.620 5.440 ;
        RECT  10.620 4.640 13.940 5.440 ;
        RECT  13.940 4.480 14.340 5.440 ;
        RECT  14.340 4.640 15.390 5.440 ;
        RECT  15.390 4.480 15.790 5.440 ;
        RECT  15.790 4.640 16.740 5.440 ;
        RECT  16.740 4.480 17.140 5.440 ;
        RECT  17.140 4.640 19.220 5.440 ;
        RECT  19.220 3.650 19.230 5.440 ;
        RECT  19.230 3.160 19.630 5.440 ;
        RECT  19.630 3.650 19.640 5.440 ;
        RECT  19.640 4.640 19.800 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        RECT  0.780 -0.400 1.180 0.560 ;
        RECT  1.180 -0.400 2.850 0.400 ;
        RECT  2.850 -0.400 3.250 0.560 ;
        RECT  3.250 -0.400 6.270 0.400 ;
        RECT  6.270 -0.400 6.670 1.440 ;
        RECT  6.670 1.200 7.890 1.440 ;
        RECT  7.890 1.200 8.290 1.600 ;
        RECT  6.670 -0.400 10.400 0.400 ;
        RECT  10.400 -0.400 10.410 0.940 ;
        RECT  10.410 -0.400 10.810 1.060 ;
        RECT  10.810 -0.400 10.820 0.940 ;
        RECT  10.820 -0.400 14.400 0.400 ;
        RECT  14.400 -0.400 14.800 0.560 ;
        RECT  14.800 -0.400 15.970 0.400 ;
        RECT  15.970 -0.400 16.950 0.560 ;
        RECT  16.950 -0.400 18.390 0.400 ;
        RECT  18.390 -0.400 18.790 0.560 ;
        RECT  18.790 -0.400 19.800 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  18.010 2.230 18.170 2.630 ;
        RECT  17.770 1.670 18.010 2.630 ;
        RECT  17.110 1.670 17.770 1.910 ;
        RECT  17.040 2.200 17.440 2.600 ;
        RECT  16.870 0.860 17.110 1.910 ;
        RECT  16.360 2.200 17.040 2.440 ;
        RECT  15.150 0.860 16.870 1.100 ;
        RECT  16.210 3.490 16.610 3.890 ;
        RECT  15.960 1.630 16.360 2.440 ;
        RECT  15.330 3.490 16.210 3.730 ;
        RECT  15.800 2.200 15.960 2.440 ;
        RECT  15.400 2.200 15.800 2.600 ;
        RECT  14.730 1.470 15.500 1.710 ;
        RECT  15.330 2.360 15.400 2.600 ;
        RECT  15.090 2.360 15.330 4.180 ;
        RECT  14.750 0.860 15.150 1.150 ;
        RECT  13.270 3.940 15.090 4.180 ;
        RECT  14.730 3.080 14.810 3.480 ;
        RECT  13.460 0.860 14.750 1.100 ;
        RECT  14.490 1.470 14.730 3.480 ;
        RECT  14.410 2.510 14.490 3.480 ;
        RECT  14.130 2.510 14.410 2.910 ;
        RECT  13.460 1.480 13.700 2.900 ;
        RECT  13.060 0.710 13.460 1.100 ;
        RECT  13.290 2.660 13.460 2.900 ;
        RECT  13.050 2.660 13.290 3.060 ;
        RECT  13.030 3.940 13.270 4.370 ;
        RECT  12.830 1.390 13.070 2.380 ;
        RECT  12.310 0.860 13.060 1.100 ;
        RECT  12.720 3.390 13.040 3.630 ;
        RECT  11.150 4.130 13.030 4.370 ;
        RECT  12.720 2.140 12.830 2.380 ;
        RECT  12.480 2.140 12.720 3.850 ;
        RECT  11.680 3.610 12.480 3.850 ;
        RECT  12.200 0.860 12.310 1.790 ;
        RECT  11.960 0.860 12.200 3.320 ;
        RECT  11.440 0.980 11.680 3.850 ;
        RECT  11.230 0.980 11.440 1.580 ;
        RECT  9.730 3.420 11.440 3.660 ;
        RECT  9.910 1.340 11.230 1.580 ;
        RECT  10.910 3.940 11.150 4.370 ;
        RECT  10.900 1.860 11.140 3.140 ;
        RECT  8.350 3.940 10.910 4.180 ;
        RECT  9.390 1.860 10.900 2.100 ;
        RECT  9.390 2.900 10.900 3.140 ;
        RECT  8.870 2.380 10.370 2.620 ;
        RECT  9.670 1.030 9.910 1.580 ;
        RECT  9.150 1.280 9.390 2.100 ;
        RECT  9.150 2.900 9.390 3.510 ;
        RECT  9.010 1.280 9.150 1.520 ;
        RECT  8.990 3.110 9.150 3.510 ;
        RECT  8.770 0.680 9.010 1.520 ;
        RECT  8.630 2.000 8.870 2.620 ;
        RECT  6.950 0.680 8.770 0.920 ;
        RECT  7.530 2.000 8.630 2.240 ;
        RECT  8.110 2.520 8.350 4.180 ;
        RECT  7.290 1.720 7.530 3.710 ;
        RECT  6.370 1.720 7.290 1.960 ;
        RECT  7.070 3.310 7.290 3.710 ;
        RECT  6.770 2.520 7.010 2.950 ;
        RECT  5.540 2.710 6.770 2.950 ;
        RECT  6.020 1.720 6.370 2.430 ;
        RECT  5.970 2.190 6.020 2.430 ;
        RECT  5.010 3.840 5.910 4.080 ;
        RECT  5.300 0.670 5.540 3.330 ;
        RECT  4.930 0.670 5.300 0.910 ;
        RECT  5.290 2.930 5.300 3.330 ;
        RECT  5.010 1.840 5.020 2.650 ;
        RECT  4.780 1.840 5.010 4.080 ;
        RECT  4.770 2.410 4.780 4.080 ;
        RECT  2.490 3.070 4.770 3.310 ;
        RECT  4.190 0.860 4.590 1.160 ;
        RECT  4.250 3.590 4.490 4.220 ;
        RECT  3.010 3.590 4.250 3.830 ;
        RECT  1.910 0.860 4.190 1.100 ;
        RECT  2.380 1.380 3.460 1.620 ;
        RECT  2.770 3.590 3.010 4.230 ;
        RECT  2.090 3.990 2.770 4.230 ;
        RECT  2.380 2.550 2.620 2.790 ;
        RECT  2.250 3.070 2.490 3.710 ;
        RECT  2.140 1.380 2.380 2.790 ;
        RECT  1.410 3.470 2.250 3.710 ;
        RECT  1.970 2.550 2.140 2.790 ;
        RECT  1.730 2.550 1.970 3.190 ;
        RECT  1.510 0.670 1.910 1.100 ;
        RECT  1.170 2.940 1.410 3.710 ;
        RECT  0.400 2.940 1.170 3.180 ;
        RECT  0.400 1.390 0.490 1.790 ;
        RECT  0.160 1.390 0.400 3.180 ;
    END
END SDFFRHQX2

MACRO SDFFRHQX1
    CLASS CORE ;
    FOREIGN SDFFRHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFRHQXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.190 2.020 3.430 2.630 ;
        RECT  3.430 2.390 3.500 2.630 ;
        RECT  3.500 2.390 3.760 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.470 1.830 1.870 2.280 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  14.410 2.910 15.070 3.260 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.120 0.710 15.290 1.110 ;
        RECT  15.290 0.710 15.520 1.480 ;
        RECT  15.520 0.790 15.530 1.480 ;
        RECT  15.920 3.780 16.050 4.180 ;
        RECT  16.040 2.950 16.050 3.210 ;
        RECT  16.050 2.950 16.100 4.180 ;
        RECT  15.530 1.240 16.100 1.480 ;
        RECT  16.100 1.240 16.340 4.180 ;
        RECT  16.340 3.130 16.350 4.180 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.880 1.740 4.510 2.100 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.180 0.860 2.640 ;
        RECT  0.860 2.180 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.650 5.440 ;
        RECT  0.650 3.770 0.890 5.440 ;
        RECT  0.890 4.640 3.290 5.440 ;
        RECT  3.290 4.110 3.530 5.440 ;
        RECT  3.530 4.640 6.300 5.440 ;
        RECT  6.300 4.140 6.310 5.440 ;
        RECT  6.310 3.940 6.710 5.440 ;
        RECT  6.710 4.140 6.720 5.440 ;
        RECT  6.720 4.640 9.530 5.440 ;
        RECT  9.530 4.480 9.930 5.440 ;
        RECT  9.930 4.640 12.450 5.440 ;
        RECT  12.450 4.480 12.850 5.440 ;
        RECT  13.740 3.070 13.900 3.310 ;
        RECT  13.900 3.070 14.140 3.770 ;
        RECT  12.850 4.640 14.700 5.440 ;
        RECT  14.140 3.530 14.700 3.770 ;
        RECT  14.700 3.530 15.100 5.440 ;
        RECT  15.100 4.640 16.500 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        RECT  0.780 -0.400 1.180 0.560 ;
        RECT  1.180 -0.400 2.850 0.400 ;
        RECT  2.850 -0.400 3.250 0.560 ;
        RECT  3.250 -0.400 6.270 0.400 ;
        RECT  6.270 -0.400 6.670 1.440 ;
        RECT  6.670 1.200 7.890 1.440 ;
        RECT  7.890 1.200 8.290 1.840 ;
        RECT  6.670 -0.400 9.200 0.400 ;
        RECT  9.200 -0.400 9.210 0.960 ;
        RECT  9.210 -0.400 9.610 1.160 ;
        RECT  9.610 -0.400 9.620 0.960 ;
        RECT  9.620 -0.400 12.140 0.400 ;
        RECT  12.140 -0.400 12.540 0.560 ;
        RECT  12.540 -0.400 13.730 0.400 ;
        RECT  13.730 -0.400 14.710 0.560 ;
        RECT  14.710 -0.400 15.910 0.400 ;
        RECT  15.910 -0.400 15.920 0.760 ;
        RECT  15.920 -0.400 16.320 0.960 ;
        RECT  16.320 -0.400 16.330 0.760 ;
        RECT  16.330 -0.400 16.500 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.660 1.760 15.820 2.000 ;
        RECT  15.340 2.400 15.580 2.810 ;
        RECT  14.100 2.400 15.340 2.640 ;
        RECT  14.420 0.860 14.660 2.000 ;
        RECT  13.050 0.860 14.420 1.100 ;
        RECT  13.380 4.050 14.340 4.290 ;
        RECT  13.700 1.380 14.100 2.640 ;
        RECT  13.440 2.050 13.700 2.640 ;
        RECT  13.380 2.400 13.440 2.640 ;
        RECT  13.140 2.400 13.380 4.290 ;
        RECT  12.700 1.470 13.250 1.710 ;
        RECT  8.430 3.940 13.140 4.180 ;
        RECT  12.500 0.860 13.050 1.150 ;
        RECT  12.700 3.210 12.860 3.450 ;
        RECT  12.460 1.470 12.700 3.450 ;
        RECT  12.040 0.860 12.500 1.100 ;
        RECT  12.340 2.550 12.460 2.950 ;
        RECT  11.800 0.860 12.040 2.350 ;
        RECT  11.110 0.860 11.800 1.110 ;
        RECT  11.790 2.110 11.800 2.350 ;
        RECT  11.550 2.110 11.790 3.660 ;
        RECT  11.110 3.420 11.550 3.660 ;
        RECT  11.270 1.590 11.520 1.830 ;
        RECT  11.030 1.590 11.270 3.140 ;
        RECT  10.870 0.860 11.110 1.310 ;
        RECT  10.550 1.590 10.750 3.650 ;
        RECT  10.510 1.060 10.550 3.650 ;
        RECT  10.310 1.060 10.510 1.830 ;
        RECT  10.350 3.410 10.510 3.650 ;
        RECT  10.030 1.060 10.310 1.300 ;
        RECT  10.030 2.300 10.230 2.700 ;
        RECT  9.790 1.580 10.030 3.660 ;
        RECT  8.810 1.580 9.790 1.820 ;
        RECT  9.050 3.420 9.790 3.660 ;
        RECT  9.270 2.170 9.510 3.140 ;
        RECT  7.530 2.170 9.270 2.410 ;
        RECT  8.570 0.680 8.810 1.820 ;
        RECT  6.950 0.680 8.570 0.920 ;
        RECT  8.190 2.690 8.430 4.180 ;
        RECT  8.030 2.690 8.190 2.930 ;
        RECT  7.290 1.720 7.530 3.710 ;
        RECT  6.180 1.720 7.290 1.960 ;
        RECT  7.070 3.310 7.290 3.710 ;
        RECT  6.770 2.550 7.010 2.950 ;
        RECT  5.540 2.710 6.770 2.950 ;
        RECT  5.940 1.720 6.180 2.400 ;
        RECT  5.010 3.790 5.910 4.030 ;
        RECT  5.530 0.670 5.540 3.250 ;
        RECT  5.300 0.670 5.530 3.330 ;
        RECT  4.930 0.670 5.300 0.910 ;
        RECT  5.290 2.930 5.300 3.330 ;
        RECT  5.010 1.800 5.020 2.650 ;
        RECT  4.780 1.800 5.010 4.030 ;
        RECT  4.770 2.370 4.780 4.030 ;
        RECT  2.490 3.070 4.770 3.310 ;
        RECT  4.190 0.860 4.590 1.200 ;
        RECT  4.250 3.590 4.490 4.070 ;
        RECT  3.010 3.590 4.250 3.830 ;
        RECT  1.910 0.860 4.190 1.100 ;
        RECT  2.380 1.380 3.460 1.620 ;
        RECT  2.770 3.590 3.010 4.230 ;
        RECT  2.090 3.990 2.770 4.230 ;
        RECT  2.380 2.550 2.620 2.790 ;
        RECT  2.250 3.070 2.490 3.710 ;
        RECT  2.140 1.380 2.380 2.790 ;
        RECT  1.410 3.470 2.250 3.710 ;
        RECT  1.970 2.550 2.140 2.790 ;
        RECT  1.730 2.550 1.970 3.190 ;
        RECT  1.670 0.670 1.910 1.100 ;
        RECT  1.510 0.670 1.670 0.910 ;
        RECT  1.170 2.940 1.410 3.710 ;
        RECT  0.400 2.940 1.170 3.180 ;
        RECT  0.400 1.260 0.490 1.660 ;
        RECT  0.160 1.260 0.400 3.180 ;
    END
END SDFFRHQX1

MACRO SDFFRXL
    CLASS CORE ;
    FOREIGN SDFFRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.820 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.150 2.020 3.500 2.640 ;
        RECT  3.500 2.020 3.550 2.650 ;
        RECT  3.550 2.390 3.760 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.440 1.830 1.780 2.350 ;
        RECT  1.780 1.950 1.860 2.350 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.800 2.950 7.060 3.210 ;
        RECT  7.060 2.950 7.470 3.200 ;
        RECT  7.470 2.950 7.770 3.190 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.880 3.670 16.040 4.070 ;
        RECT  16.040 3.510 16.380 4.070 ;
        RECT  15.990 0.730 16.390 1.100 ;
        RECT  16.380 3.520 16.730 3.760 ;
        RECT  16.390 0.860 16.730 1.100 ;
        RECT  16.730 0.860 16.970 3.760 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.250 1.390 17.270 1.790 ;
        RECT  17.270 1.390 17.360 1.820 ;
        RECT  17.250 2.980 17.370 3.380 ;
        RECT  17.360 1.390 17.370 2.090 ;
        RECT  17.370 1.390 17.610 3.380 ;
        RECT  17.610 1.830 17.620 2.090 ;
        RECT  17.610 2.980 17.650 3.380 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.000 1.700 4.510 2.120 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 0.870 3.210 ;
        RECT  0.710 2.070 0.870 2.470 ;
        RECT  0.870 2.070 1.110 3.210 ;
        RECT  1.110 2.950 1.120 3.210 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.380 5.440 ;
        RECT  0.380 4.480 2.020 5.440 ;
        RECT  2.020 4.640 3.350 5.440 ;
        RECT  3.350 4.310 3.360 5.440 ;
        RECT  3.360 4.190 3.760 5.440 ;
        RECT  3.760 4.310 3.770 5.440 ;
        RECT  3.770 4.640 6.730 5.440 ;
        RECT  6.730 4.480 7.130 5.440 ;
        RECT  7.130 4.640 10.300 5.440 ;
        RECT  10.300 4.110 11.280 5.440 ;
        RECT  11.280 4.640 13.150 5.440 ;
        RECT  13.150 4.170 13.160 5.440 ;
        RECT  13.160 3.970 13.560 5.440 ;
        RECT  13.560 4.170 13.570 5.440 ;
        RECT  13.570 4.640 15.110 5.440 ;
        RECT  15.110 3.860 15.120 5.440 ;
        RECT  15.120 3.660 15.520 5.440 ;
        RECT  15.520 3.860 15.530 5.440 ;
        RECT  15.530 4.640 17.140 5.440 ;
        RECT  17.140 4.480 17.540 5.440 ;
        RECT  17.540 4.640 17.820 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        RECT  0.900 -0.400 1.300 0.560 ;
        RECT  1.300 -0.400 2.970 0.400 ;
        RECT  2.970 -0.400 3.370 0.560 ;
        RECT  3.370 -0.400 6.610 0.400 ;
        RECT  6.610 -0.400 6.620 0.730 ;
        RECT  6.620 -0.400 7.020 0.850 ;
        RECT  7.020 -0.400 7.030 0.730 ;
        RECT  7.030 -0.400 8.870 0.400 ;
        RECT  8.870 -0.400 9.130 1.530 ;
        RECT  9.130 1.290 10.640 1.530 ;
        RECT  10.640 1.270 10.650 1.600 ;
        RECT  10.650 1.270 11.050 1.820 ;
        RECT  11.050 1.270 11.060 1.600 ;
        RECT  9.130 -0.400 13.330 0.400 ;
        RECT  13.330 -0.400 13.340 1.090 ;
        RECT  13.340 -0.400 13.740 1.290 ;
        RECT  13.740 -0.400 13.750 1.090 ;
        RECT  13.750 -0.400 15.090 0.400 ;
        RECT  15.090 -0.400 15.100 0.890 ;
        RECT  15.100 -0.400 15.500 1.090 ;
        RECT  15.500 -0.400 15.510 0.890 ;
        RECT  15.510 -0.400 17.050 0.400 ;
        RECT  17.050 -0.400 17.450 0.560 ;
        RECT  17.450 -0.400 17.820 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.210 1.470 16.450 3.180 ;
        RECT  15.990 1.470 16.210 1.710 ;
        RECT  15.910 2.780 16.210 3.180 ;
        RECT  14.980 1.970 15.740 2.370 ;
        RECT  14.740 1.590 14.980 3.270 ;
        RECT  14.620 1.590 14.740 1.830 ;
        RECT  14.300 3.030 14.740 3.270 ;
        RECT  14.220 1.030 14.620 1.830 ;
        RECT  14.060 2.170 14.460 2.570 ;
        RECT  14.060 3.030 14.300 4.010 ;
        RECT  13.460 1.590 14.220 1.830 ;
        RECT  12.780 2.330 14.060 2.570 ;
        RECT  13.900 3.610 14.060 4.010 ;
        RECT  13.060 1.590 13.460 1.990 ;
        RECT  12.780 3.730 12.820 4.130 ;
        RECT  12.770 2.330 12.780 4.130 ;
        RECT  12.530 1.180 12.770 4.130 ;
        RECT  12.400 1.180 12.530 1.420 ;
        RECT  12.420 3.730 12.530 4.130 ;
        RECT  12.000 1.020 12.400 1.420 ;
        RECT  12.140 2.380 12.220 2.780 ;
        RECT  11.900 2.380 12.140 3.830 ;
        RECT  11.620 1.740 12.100 1.980 ;
        RECT  10.420 3.590 11.900 3.830 ;
        RECT  11.380 0.670 11.620 3.310 ;
        RECT  9.410 0.670 11.380 0.910 ;
        RECT  10.700 3.070 11.380 3.310 ;
        RECT  9.770 2.160 11.100 2.560 ;
        RECT  10.180 2.880 10.420 3.830 ;
        RECT  9.710 3.590 10.180 3.830 ;
        RECT  9.530 1.820 9.770 3.140 ;
        RECT  9.470 3.590 9.710 4.290 ;
        RECT  8.590 1.820 9.530 2.060 ;
        RECT  9.080 2.900 9.530 3.140 ;
        RECT  7.660 4.050 9.470 4.290 ;
        RECT  8.340 2.340 9.250 2.580 ;
        RECT  8.840 2.900 9.080 3.770 ;
        RECT  8.680 3.530 8.840 3.770 ;
        RECT  8.350 1.110 8.590 2.060 ;
        RECT  8.220 1.110 8.350 1.890 ;
        RECT  8.100 2.340 8.340 3.770 ;
        RECT  6.490 1.650 8.220 1.890 ;
        RECT  8.070 2.340 8.100 2.580 ;
        RECT  7.940 3.530 8.100 3.770 ;
        RECT  7.670 2.170 8.070 2.580 ;
        RECT  7.540 0.770 7.940 1.010 ;
        RECT  7.420 3.940 7.660 4.290 ;
        RECT  7.300 0.770 7.540 1.370 ;
        RECT  6.450 3.940 7.420 4.180 ;
        RECT  5.970 1.130 7.300 1.370 ;
        RECT  6.250 1.650 6.490 2.080 ;
        RECT  5.690 3.940 6.450 4.320 ;
        RECT  5.970 2.360 6.210 3.650 ;
        RECT  5.730 1.130 5.970 2.600 ;
        RECT  5.530 1.130 5.730 1.370 ;
        RECT  5.450 2.880 5.690 4.320 ;
        RECT  5.130 0.930 5.530 1.370 ;
        RECT  5.210 1.680 5.450 3.120 ;
        RECT  4.280 4.080 5.450 4.320 ;
        RECT  4.830 1.680 5.210 2.080 ;
        RECT  4.930 3.400 5.170 3.800 ;
        RECT  4.690 3.150 4.930 3.800 ;
        RECT  4.310 0.860 4.710 1.330 ;
        RECT  2.390 3.150 4.690 3.390 ;
        RECT  2.220 0.860 4.310 1.100 ;
        RECT  4.040 3.670 4.280 4.320 ;
        RECT  3.060 3.670 4.040 3.910 ;
        RECT  2.380 1.380 3.670 1.620 ;
        RECT  2.820 3.670 3.060 3.990 ;
        RECT  2.380 2.470 2.830 2.870 ;
        RECT  0.500 3.750 2.820 3.990 ;
        RECT  2.140 1.380 2.380 2.870 ;
        RECT  1.980 0.670 2.220 1.100 ;
        RECT  2.050 2.630 2.140 2.870 ;
        RECT  1.810 2.630 2.050 3.470 ;
        RECT  1.630 0.670 1.980 0.910 ;
        RECT  1.650 3.070 1.810 3.470 ;
        RECT  0.410 1.300 0.570 1.700 ;
        RECT  0.410 2.930 0.500 3.990 ;
        RECT  0.260 1.300 0.410 3.990 ;
        RECT  0.170 1.300 0.260 3.360 ;
    END
END SDFFRXL

MACRO SDFFRX4
    CLASS CORE ;
    FOREIGN SDFFRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFRXL ;
    SIZE 23.100 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.650 2.160 3.170 2.660 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.270 1.570 1.530 ;
        RECT  1.570 1.270 1.780 2.340 ;
        RECT  1.780 1.290 1.810 2.340 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.310 2.610 7.320 3.050 ;
        RECT  7.320 2.610 7.720 3.210 ;
        RECT  7.720 2.610 7.730 3.050 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  20.420 2.750 20.550 3.150 ;
        RECT  20.550 1.170 20.570 3.150 ;
        RECT  20.570 1.170 20.950 3.220 ;
        RECT  20.950 1.820 21.010 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.880 2.720 21.890 3.160 ;
        RECT  21.890 1.170 22.290 3.160 ;
        RECT  22.290 1.260 22.330 3.160 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.020 1.620 4.510 2.100 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.700 2.150 0.710 2.570 ;
        RECT  0.710 2.150 0.860 2.640 ;
        RECT  0.860 2.150 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.200 5.440 ;
        RECT  0.200 4.480 0.600 5.440 ;
        RECT  0.600 4.640 2.380 5.440 ;
        RECT  2.380 3.940 3.360 5.440 ;
        RECT  3.360 4.640 6.880 5.440 ;
        RECT  6.880 4.480 7.280 5.440 ;
        RECT  7.280 4.640 10.470 5.440 ;
        RECT  10.470 4.180 12.010 5.440 ;
        RECT  12.010 4.640 14.550 5.440 ;
        RECT  14.550 4.290 14.560 5.440 ;
        RECT  14.560 4.090 14.960 5.440 ;
        RECT  14.960 4.290 14.970 5.440 ;
        RECT  14.970 4.640 15.870 5.440 ;
        RECT  15.870 4.280 15.880 5.440 ;
        RECT  15.880 4.080 16.280 5.440 ;
        RECT  16.280 4.280 16.290 5.440 ;
        RECT  16.290 4.640 18.350 5.440 ;
        RECT  18.350 3.450 18.360 5.440 ;
        RECT  18.360 2.960 18.760 5.440 ;
        RECT  18.760 3.450 18.770 5.440 ;
        RECT  18.770 4.640 19.740 5.440 ;
        RECT  19.740 4.210 19.750 5.440 ;
        RECT  19.750 4.010 20.150 5.440 ;
        RECT  20.150 4.210 20.160 5.440 ;
        RECT  20.160 4.640 21.130 5.440 ;
        RECT  21.130 4.210 21.140 5.440 ;
        RECT  21.140 4.010 21.540 5.440 ;
        RECT  21.540 4.210 21.550 5.440 ;
        RECT  21.550 4.640 22.520 5.440 ;
        RECT  22.520 4.210 22.530 5.440 ;
        RECT  22.530 4.010 22.930 5.440 ;
        RECT  22.930 4.210 22.940 5.440 ;
        RECT  22.940 4.640 23.100 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.920 0.400 ;
        RECT  0.920 -0.400 1.320 0.560 ;
        RECT  1.320 -0.400 3.010 0.400 ;
        RECT  3.010 -0.400 3.410 0.560 ;
        RECT  3.410 -0.400 7.670 0.400 ;
        RECT  7.670 -0.400 8.650 1.290 ;
        RECT  8.650 -0.400 9.580 0.400 ;
        RECT  9.580 -0.400 9.590 0.890 ;
        RECT  9.590 -0.400 9.990 1.090 ;
        RECT  9.990 -0.400 10.000 0.890 ;
        RECT  10.000 -0.400 11.290 0.400 ;
        RECT  11.290 -0.400 11.300 1.120 ;
        RECT  11.300 -0.400 11.700 1.320 ;
        RECT  11.700 -0.400 11.710 1.120 ;
        RECT  11.710 -0.400 13.880 0.400 ;
        RECT  13.880 -0.400 13.890 0.890 ;
        RECT  13.890 -0.400 14.290 1.090 ;
        RECT  14.290 -0.400 14.300 0.890 ;
        RECT  14.300 -0.400 16.360 0.400 ;
        RECT  16.360 -0.400 17.340 1.010 ;
        RECT  17.340 -0.400 18.380 0.400 ;
        RECT  18.380 -0.400 18.390 1.130 ;
        RECT  18.390 -0.400 18.790 1.620 ;
        RECT  18.790 -0.400 18.800 1.130 ;
        RECT  18.800 -0.400 19.900 0.400 ;
        RECT  19.900 -0.400 19.910 0.680 ;
        RECT  19.910 -0.400 20.310 0.880 ;
        RECT  20.310 -0.400 20.320 0.680 ;
        RECT  20.320 -0.400 21.210 0.400 ;
        RECT  21.210 -0.400 21.220 0.690 ;
        RECT  21.220 -0.400 21.620 0.890 ;
        RECT  21.620 -0.400 21.630 0.690 ;
        RECT  21.630 -0.400 22.500 0.400 ;
        RECT  22.500 -0.400 22.510 0.690 ;
        RECT  22.510 -0.400 22.910 0.890 ;
        RECT  22.910 -0.400 22.920 0.690 ;
        RECT  22.920 -0.400 23.100 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  22.600 2.180 22.840 3.730 ;
        RECT  20.140 3.490 22.600 3.730 ;
        RECT  19.900 1.550 20.140 3.730 ;
        RECT  19.590 1.550 19.900 1.790 ;
        RECT  19.080 3.270 19.900 3.670 ;
        RECT  18.070 2.070 19.620 2.470 ;
        RECT  19.190 1.390 19.590 1.790 ;
        RECT  17.830 0.660 18.070 3.490 ;
        RECT  17.670 0.660 17.830 1.640 ;
        RECT  17.630 3.250 17.830 3.490 ;
        RECT  16.070 1.390 17.670 1.630 ;
        RECT  17.160 3.250 17.630 3.790 ;
        RECT  16.920 2.200 17.320 2.600 ;
        RECT  15.600 3.550 17.160 3.790 ;
        RECT  15.700 2.200 16.920 2.530 ;
        RECT  15.820 1.160 16.070 1.630 ;
        RECT  15.670 1.160 15.820 1.400 ;
        RECT  15.540 2.130 15.700 2.530 ;
        RECT  15.360 3.550 15.600 4.350 ;
        RECT  15.300 1.820 15.540 3.270 ;
        RECT  15.100 1.820 15.300 2.060 ;
        RECT  14.910 3.030 15.300 3.270 ;
        RECT  14.860 0.690 15.100 2.060 ;
        RECT  14.780 2.340 15.020 2.740 ;
        RECT  14.670 3.030 14.910 3.590 ;
        RECT  14.630 0.690 14.860 1.620 ;
        RECT  14.580 2.340 14.780 2.580 ;
        RECT  13.680 3.350 14.670 3.590 ;
        RECT  13.400 1.380 14.630 1.620 ;
        RECT  14.340 1.900 14.580 2.580 ;
        RECT  12.680 1.900 14.340 2.140 ;
        RECT  12.890 2.690 13.930 2.930 ;
        RECT  13.280 3.350 13.680 3.860 ;
        RECT  13.160 1.190 13.400 1.620 ;
        RECT  12.520 1.190 13.160 1.430 ;
        RECT  12.650 2.690 12.890 3.900 ;
        RECT  12.600 1.730 12.680 2.140 ;
        RECT  11.010 3.660 12.650 3.900 ;
        RECT  12.360 1.710 12.600 2.140 ;
        RECT  12.120 1.710 12.360 3.160 ;
        RECT  10.740 1.710 12.120 1.950 ;
        RECT  11.530 2.920 12.120 3.160 ;
        RECT  10.180 2.250 11.840 2.490 ;
        RECT  11.290 2.920 11.530 3.380 ;
        RECT  10.770 2.770 11.010 3.900 ;
        RECT  10.610 2.770 10.770 3.540 ;
        RECT  10.500 0.670 10.740 1.950 ;
        RECT  10.110 3.300 10.610 3.540 ;
        RECT  10.280 0.670 10.500 0.910 ;
        RECT  9.940 1.570 10.180 3.020 ;
        RECT  9.870 3.300 10.110 4.270 ;
        RECT  6.840 1.570 9.940 1.810 ;
        RECT  9.590 2.780 9.940 3.020 ;
        RECT  7.810 4.030 9.870 4.270 ;
        RECT  8.330 2.150 9.660 2.390 ;
        RECT  9.350 2.780 9.590 3.690 ;
        RECT  9.190 3.450 9.350 3.690 ;
        RECT  8.330 3.510 8.660 3.750 ;
        RECT  8.090 2.090 8.330 3.750 ;
        RECT  8.080 2.090 8.090 2.390 ;
        RECT  7.640 2.090 8.080 2.330 ;
        RECT  7.570 3.940 7.810 4.270 ;
        RECT  6.470 3.940 7.570 4.180 ;
        RECT  5.810 0.770 7.400 1.010 ;
        RECT  6.600 1.570 6.840 2.690 ;
        RECT  6.440 2.290 6.600 2.690 ;
        RECT  6.230 3.940 6.470 4.350 ;
        RECT  5.290 4.110 6.230 4.350 ;
        RECT  5.570 0.770 5.810 3.830 ;
        RECT  5.380 1.090 5.570 1.490 ;
        RECT  5.050 1.880 5.290 4.350 ;
        RECT  4.840 1.880 5.050 2.280 ;
        RECT  4.110 4.110 5.050 4.350 ;
        RECT  4.420 0.860 4.820 1.350 ;
        RECT  4.530 2.860 4.770 3.830 ;
        RECT  3.600 2.860 4.530 3.100 ;
        RECT  2.730 0.860 4.420 1.100 ;
        RECT  3.870 3.420 4.110 4.350 ;
        RECT  0.570 3.420 3.870 3.660 ;
        RECT  3.310 1.380 3.710 1.780 ;
        RECT  2.380 1.540 3.310 1.780 ;
        RECT  2.490 0.670 2.730 1.100 ;
        RECT  1.650 0.670 2.490 0.910 ;
        RECT  2.140 1.430 2.380 3.090 ;
        RECT  1.650 2.850 2.140 3.090 ;
        RECT  0.410 1.190 0.570 1.590 ;
        RECT  0.410 3.010 0.570 3.660 ;
        RECT  0.330 1.190 0.410 3.660 ;
        RECT  0.170 1.190 0.330 3.410 ;
    END
END SDFFRX4

MACRO SDFFRX2
    CLASS CORE ;
    FOREIGN SDFFRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFRXL ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.770 2.020 2.840 2.640 ;
        RECT  2.840 2.020 3.100 2.650 ;
        RECT  3.100 2.020 3.170 2.420 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 1.280 1.520 2.300 ;
        RECT  1.520 1.270 1.720 2.300 ;
        RECT  1.720 1.270 1.780 1.530 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.800 2.950 6.810 3.210 ;
        RECT  6.810 2.710 7.060 3.210 ;
        RECT  7.060 2.710 7.560 3.110 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.040 2.920 17.120 3.320 ;
        RECT  17.120 2.610 17.130 3.320 ;
        RECT  17.040 0.730 17.130 1.710 ;
        RECT  17.130 0.730 17.370 3.320 ;
        RECT  17.370 2.390 17.440 3.320 ;
        RECT  17.370 0.730 17.440 1.710 ;
        RECT  17.440 2.390 17.620 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.570 0.730 18.680 1.830 ;
        RECT  18.570 3.170 18.690 4.150 ;
        RECT  18.680 0.730 18.690 2.090 ;
        RECT  18.690 0.730 18.930 4.150 ;
        RECT  18.930 0.730 18.940 2.090 ;
        RECT  18.930 3.170 18.970 4.150 ;
        RECT  18.940 0.730 18.970 1.960 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.940 1.510 4.420 2.100 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.060 0.770 2.460 ;
        RECT  0.770 1.820 1.130 2.470 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.260 5.440 ;
        RECT  0.260 4.480 0.660 5.440 ;
        RECT  0.660 4.640 3.670 5.440 ;
        RECT  3.670 4.090 4.070 5.440 ;
        RECT  4.070 4.640 6.650 5.440 ;
        RECT  6.650 4.480 7.050 5.440 ;
        RECT  7.050 4.640 9.950 5.440 ;
        RECT  9.950 4.170 11.490 5.440 ;
        RECT  11.490 4.640 13.510 5.440 ;
        RECT  13.510 4.110 13.520 5.440 ;
        RECT  13.520 3.910 13.920 5.440 ;
        RECT  13.920 4.110 13.930 5.440 ;
        RECT  13.930 4.640 15.470 5.440 ;
        RECT  15.470 3.500 15.480 5.440 ;
        RECT  15.480 3.300 15.880 5.440 ;
        RECT  15.880 3.500 15.890 5.440 ;
        RECT  15.890 4.640 17.800 5.440 ;
        RECT  17.800 4.320 17.810 5.440 ;
        RECT  17.810 4.120 18.210 5.440 ;
        RECT  18.210 4.320 18.220 5.440 ;
        RECT  18.220 4.640 19.140 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 2.910 0.400 ;
        RECT  2.910 -0.400 3.310 0.560 ;
        RECT  3.310 -0.400 7.510 0.400 ;
        RECT  7.510 -0.400 7.910 1.310 ;
        RECT  7.910 -0.400 9.000 0.400 ;
        RECT  9.000 -0.400 9.010 0.640 ;
        RECT  9.010 -0.400 9.410 0.930 ;
        RECT  9.410 -0.400 9.420 0.640 ;
        RECT  9.420 -0.400 10.700 0.400 ;
        RECT  10.700 -0.400 10.710 1.020 ;
        RECT  10.710 -0.400 11.110 1.140 ;
        RECT  11.110 -0.400 11.120 1.020 ;
        RECT  11.120 -0.400 13.790 0.400 ;
        RECT  13.790 -0.400 14.190 0.560 ;
        RECT  14.190 -0.400 15.360 0.400 ;
        RECT  15.360 -0.400 15.370 1.100 ;
        RECT  15.370 -0.400 15.770 1.300 ;
        RECT  15.770 -0.400 15.780 1.100 ;
        RECT  15.780 -0.400 17.800 0.400 ;
        RECT  17.800 -0.400 17.810 1.200 ;
        RECT  17.810 -0.400 18.210 1.690 ;
        RECT  18.210 -0.400 18.220 1.200 ;
        RECT  18.220 -0.400 19.140 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  18.290 2.200 18.320 2.600 ;
        RECT  18.050 2.200 18.290 3.840 ;
        RECT  16.760 3.600 18.050 3.840 ;
        RECT  16.520 1.080 16.760 3.840 ;
        RECT  16.190 1.080 16.520 1.480 ;
        RECT  16.300 2.920 16.520 3.320 ;
        RECT  15.290 1.950 16.240 2.350 ;
        RECT  15.050 1.580 15.290 3.020 ;
        RECT  15.010 1.580 15.050 1.820 ;
        RECT  14.660 2.780 15.050 3.020 ;
        RECT  14.610 0.940 15.010 1.820 ;
        RECT  14.370 2.100 14.770 2.500 ;
        RECT  14.420 2.780 14.660 3.900 ;
        RECT  13.740 1.580 14.610 1.820 ;
        RECT  14.260 2.920 14.420 3.900 ;
        RECT  13.060 2.260 14.370 2.500 ;
        RECT  13.340 1.580 13.740 1.980 ;
        RECT  12.820 1.260 13.060 3.490 ;
        RECT  12.390 1.260 12.820 1.500 ;
        RECT  12.700 3.250 12.820 3.490 ;
        RECT  12.460 3.250 12.700 3.650 ;
        RECT  12.120 2.610 12.540 2.850 ;
        RECT  11.990 1.100 12.390 1.500 ;
        RECT  11.600 1.890 12.130 2.130 ;
        RECT  11.880 2.610 12.120 3.890 ;
        RECT  10.260 3.650 11.880 3.890 ;
        RECT  11.360 1.420 11.600 3.350 ;
        RECT  10.230 1.420 11.360 1.710 ;
        RECT  10.540 3.110 11.360 3.350 ;
        RECT  10.840 1.990 11.080 2.710 ;
        RECT  9.490 1.990 10.840 2.230 ;
        RECT  10.260 2.510 10.440 2.750 ;
        RECT  10.020 2.510 10.260 3.890 ;
        RECT  10.100 1.310 10.230 1.710 ;
        RECT  10.090 0.880 10.100 1.710 ;
        RECT  9.830 0.670 10.090 1.710 ;
        RECT  9.580 3.650 10.020 3.890 ;
        RECT  9.690 0.670 9.830 0.910 ;
        RECT  9.340 3.650 9.580 4.310 ;
        RECT  9.250 1.590 9.490 3.190 ;
        RECT  7.570 4.070 9.340 4.310 ;
        RECT  8.830 1.590 9.250 1.830 ;
        RECT  9.020 2.950 9.250 3.190 ;
        RECT  8.780 2.950 9.020 3.790 ;
        RECT  8.730 2.110 8.970 2.510 ;
        RECT  8.430 1.270 8.830 1.830 ;
        RECT  8.620 3.390 8.780 3.790 ;
        RECT  8.090 2.110 8.730 2.350 ;
        RECT  6.570 1.590 8.430 1.830 ;
        RECT  7.850 2.110 8.090 3.790 ;
        RECT  7.550 2.110 7.850 2.350 ;
        RECT  7.330 3.940 7.570 4.310 ;
        RECT  6.350 3.940 7.330 4.180 ;
        RECT  6.830 0.670 7.230 1.090 ;
        RECT  5.830 0.670 6.830 0.910 ;
        RECT  6.330 1.590 6.570 2.270 ;
        RECT  6.110 3.940 6.350 4.250 ;
        RECT  6.170 1.870 6.330 2.270 ;
        RECT  5.310 4.010 6.110 4.250 ;
        RECT  5.590 0.670 5.830 3.490 ;
        RECT  5.130 0.800 5.590 1.200 ;
        RECT  5.070 1.500 5.310 4.250 ;
        RECT  4.830 1.500 5.070 1.900 ;
        RECT  4.650 4.010 5.070 4.250 ;
        RECT  4.550 2.770 4.790 3.170 ;
        RECT  4.250 0.860 4.650 1.220 ;
        RECT  4.410 3.450 4.650 4.250 ;
        RECT  2.770 2.930 4.550 3.170 ;
        RECT  3.290 3.450 4.410 3.690 ;
        RECT  2.570 0.860 4.250 1.100 ;
        RECT  2.380 1.380 3.610 1.620 ;
        RECT  3.050 3.450 3.290 4.220 ;
        RECT  1.510 3.980 3.050 4.220 ;
        RECT  2.530 2.930 2.770 3.330 ;
        RECT  2.330 0.670 2.570 1.100 ;
        RECT  2.250 1.380 2.380 2.050 ;
        RECT  1.570 0.670 2.330 0.910 ;
        RECT  2.140 1.380 2.250 3.700 ;
        RECT  2.010 1.810 2.140 3.700 ;
        RECT  1.790 2.810 2.010 3.700 ;
        RECT  1.270 3.080 1.510 4.220 ;
        RECT  0.570 3.080 1.270 3.320 ;
        RECT  0.400 2.920 0.570 3.320 ;
        RECT  0.400 1.310 0.490 1.710 ;
        RECT  0.160 1.310 0.400 3.320 ;
    END
END SDFFRX2

MACRO SDFFRX1
    CLASS CORE ;
    FOREIGN SDFFRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFRXL ;
    SIZE 17.820 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.150 2.020 3.500 2.640 ;
        RECT  3.500 2.020 3.550 2.650 ;
        RECT  3.550 2.390 3.760 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.440 1.830 1.780 2.350 ;
        RECT  1.780 1.950 1.860 2.350 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.800 2.950 7.060 3.210 ;
        RECT  7.060 2.950 7.470 3.200 ;
        RECT  7.470 2.950 7.770 3.190 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.900 3.670 16.040 4.070 ;
        RECT  15.840 0.710 16.250 1.100 ;
        RECT  16.040 3.510 16.380 4.070 ;
        RECT  16.380 3.520 16.730 3.760 ;
        RECT  16.250 0.860 16.730 1.100 ;
        RECT  16.730 0.860 16.970 3.760 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.250 1.320 17.270 1.720 ;
        RECT  17.270 1.320 17.360 1.820 ;
        RECT  17.250 2.980 17.370 3.380 ;
        RECT  17.360 1.320 17.370 2.090 ;
        RECT  17.370 1.320 17.610 3.380 ;
        RECT  17.610 1.320 17.620 2.090 ;
        RECT  17.610 2.980 17.650 3.380 ;
        RECT  17.620 1.320 17.650 1.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.940 1.640 3.950 2.100 ;
        RECT  3.950 1.610 4.410 2.100 ;
        RECT  4.410 1.640 4.420 2.100 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 0.870 3.210 ;
        RECT  0.710 2.070 0.870 2.470 ;
        RECT  0.870 2.070 1.110 3.210 ;
        RECT  1.110 2.950 1.120 3.210 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.980 5.440 ;
        RECT  0.980 4.480 2.020 5.440 ;
        RECT  2.020 4.640 3.350 5.440 ;
        RECT  3.350 4.310 3.360 5.440 ;
        RECT  3.360 4.190 3.760 5.440 ;
        RECT  3.760 4.310 3.770 5.440 ;
        RECT  3.770 4.640 6.730 5.440 ;
        RECT  6.730 4.480 7.130 5.440 ;
        RECT  7.130 4.640 10.300 5.440 ;
        RECT  10.300 4.110 11.280 5.440 ;
        RECT  11.280 4.640 13.150 5.440 ;
        RECT  13.150 4.170 13.160 5.440 ;
        RECT  13.160 3.970 13.560 5.440 ;
        RECT  13.560 4.170 13.570 5.440 ;
        RECT  13.570 4.640 15.130 5.440 ;
        RECT  15.130 3.860 15.140 5.440 ;
        RECT  15.140 3.660 15.540 5.440 ;
        RECT  15.540 3.860 15.550 5.440 ;
        RECT  15.550 4.640 16.650 5.440 ;
        RECT  16.650 4.480 17.050 5.440 ;
        RECT  17.050 4.640 17.820 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 2.910 0.400 ;
        RECT  2.910 -0.400 3.310 0.560 ;
        RECT  3.310 -0.400 6.610 0.400 ;
        RECT  6.610 -0.400 6.620 0.730 ;
        RECT  6.620 -0.400 7.020 0.850 ;
        RECT  7.020 -0.400 7.030 0.730 ;
        RECT  7.030 -0.400 8.870 0.400 ;
        RECT  8.870 -0.400 9.130 1.530 ;
        RECT  9.130 1.290 10.640 1.530 ;
        RECT  10.640 1.270 10.650 1.600 ;
        RECT  10.650 1.270 11.050 1.820 ;
        RECT  11.050 1.270 11.060 1.600 ;
        RECT  9.130 -0.400 13.340 0.400 ;
        RECT  13.340 -0.400 13.740 1.270 ;
        RECT  13.740 -0.400 15.080 0.400 ;
        RECT  15.080 -0.400 15.090 0.690 ;
        RECT  15.090 -0.400 15.490 0.890 ;
        RECT  15.490 -0.400 15.500 0.690 ;
        RECT  15.500 -0.400 17.140 0.400 ;
        RECT  17.140 -0.400 17.540 0.560 ;
        RECT  17.540 -0.400 17.820 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.210 1.450 16.450 3.180 ;
        RECT  15.910 1.450 16.210 1.690 ;
        RECT  15.910 2.780 16.210 3.180 ;
        RECT  14.980 1.970 15.740 2.370 ;
        RECT  14.740 1.590 14.980 3.270 ;
        RECT  14.650 1.590 14.740 1.830 ;
        RECT  14.320 3.030 14.740 3.270 ;
        RECT  14.250 0.880 14.650 1.830 ;
        RECT  14.060 2.150 14.460 2.550 ;
        RECT  13.920 3.030 14.320 3.640 ;
        RECT  13.460 1.590 14.250 1.830 ;
        RECT  12.780 2.270 14.060 2.510 ;
        RECT  13.060 1.590 13.460 1.990 ;
        RECT  12.780 3.730 12.820 4.130 ;
        RECT  12.770 2.270 12.780 4.130 ;
        RECT  12.530 1.180 12.770 4.130 ;
        RECT  12.400 1.180 12.530 1.420 ;
        RECT  12.420 3.730 12.530 4.130 ;
        RECT  12.000 1.020 12.400 1.420 ;
        RECT  12.140 2.490 12.220 2.890 ;
        RECT  11.900 2.490 12.140 3.830 ;
        RECT  11.620 1.850 12.100 2.090 ;
        RECT  10.420 3.590 11.900 3.830 ;
        RECT  11.380 0.670 11.620 3.310 ;
        RECT  9.410 0.670 11.380 0.910 ;
        RECT  10.700 3.070 11.380 3.310 ;
        RECT  9.770 2.160 11.100 2.560 ;
        RECT  10.180 2.880 10.420 3.830 ;
        RECT  9.710 3.590 10.180 3.830 ;
        RECT  9.530 1.820 9.770 3.140 ;
        RECT  9.470 3.590 9.710 4.290 ;
        RECT  8.590 1.820 9.530 2.060 ;
        RECT  9.080 2.900 9.530 3.140 ;
        RECT  7.660 4.050 9.470 4.290 ;
        RECT  8.340 2.340 9.250 2.580 ;
        RECT  8.840 2.900 9.080 3.770 ;
        RECT  8.680 3.530 8.840 3.770 ;
        RECT  8.350 1.110 8.590 2.060 ;
        RECT  8.220 1.110 8.350 1.890 ;
        RECT  8.100 2.340 8.340 3.770 ;
        RECT  6.490 1.650 8.220 1.890 ;
        RECT  8.070 2.340 8.100 2.580 ;
        RECT  7.940 3.530 8.100 3.770 ;
        RECT  7.670 2.170 8.070 2.580 ;
        RECT  7.540 0.770 7.940 1.010 ;
        RECT  7.420 3.940 7.660 4.290 ;
        RECT  7.300 0.770 7.540 1.370 ;
        RECT  6.450 3.940 7.420 4.180 ;
        RECT  5.970 1.130 7.300 1.370 ;
        RECT  6.250 1.650 6.490 2.080 ;
        RECT  5.690 3.940 6.450 4.320 ;
        RECT  5.970 2.360 6.210 3.650 ;
        RECT  5.730 1.130 5.970 2.600 ;
        RECT  5.530 1.130 5.730 1.370 ;
        RECT  5.450 2.880 5.690 4.320 ;
        RECT  5.130 0.930 5.530 1.370 ;
        RECT  5.210 1.680 5.450 3.120 ;
        RECT  4.280 4.080 5.450 4.320 ;
        RECT  4.830 1.680 5.210 2.080 ;
        RECT  4.930 3.400 5.170 3.800 ;
        RECT  4.690 3.150 4.930 3.800 ;
        RECT  2.390 3.150 4.690 3.390 ;
        RECT  4.250 0.860 4.650 1.330 ;
        RECT  4.040 3.670 4.280 4.320 ;
        RECT  2.160 0.860 4.250 1.100 ;
        RECT  2.620 3.670 4.040 3.910 ;
        RECT  2.380 1.380 3.610 1.620 ;
        RECT  2.380 2.470 2.830 2.870 ;
        RECT  2.380 3.670 2.620 3.990 ;
        RECT  2.140 1.380 2.380 2.870 ;
        RECT  0.490 3.750 2.380 3.990 ;
        RECT  1.920 0.670 2.160 1.100 ;
        RECT  2.050 2.630 2.140 2.870 ;
        RECT  1.810 2.630 2.050 3.470 ;
        RECT  1.570 0.670 1.920 0.910 ;
        RECT  1.650 3.070 1.810 3.470 ;
        RECT  0.410 1.300 0.570 1.700 ;
        RECT  0.410 2.930 0.490 3.990 ;
        RECT  0.250 1.300 0.410 3.990 ;
        RECT  0.170 1.300 0.250 3.360 ;
    END
END SDFFRX1

MACRO SDFFNSRXL
    CLASS CORE ;
    FOREIGN SDFFNSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.920 3.940 7.320 4.370 ;
        RECT  7.320 3.940 8.530 4.180 ;
        RECT  8.530 3.940 8.770 4.360 ;
        RECT  8.770 4.080 8.790 4.360 ;
        RECT  8.790 4.120 10.700 4.360 ;
        RECT  10.700 4.120 10.940 4.370 ;
        RECT  10.940 4.130 14.550 4.370 ;
        RECT  14.550 3.930 14.970 4.370 ;
        RECT  14.970 4.070 14.980 4.370 ;
        RECT  14.980 4.080 15.010 4.370 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.950 2.850 3.210 ;
        RECT  2.850 2.180 3.090 3.210 ;
        RECT  3.090 2.950 3.100 3.210 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.950 0.210 3.210 ;
        RECT  0.210 2.560 0.460 3.210 ;
        RECT  0.460 2.560 0.530 3.200 ;
        RECT  0.530 2.560 0.610 2.960 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.120 1.270 8.380 1.530 ;
        RECT  8.380 1.280 8.430 1.530 ;
        RECT  8.430 1.280 8.670 1.890 ;
        RECT  8.670 1.650 8.710 1.890 ;
        RECT  8.710 1.650 8.950 2.110 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.810 1.390 17.210 1.790 ;
        RECT  16.930 2.960 17.360 3.200 ;
        RECT  17.360 2.950 17.530 3.210 ;
        RECT  17.210 1.550 17.530 1.790 ;
        RECT  17.530 1.550 17.620 3.210 ;
        RECT  17.620 1.550 17.770 3.200 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.570 2.940 18.690 3.340 ;
        RECT  18.680 2.390 18.690 2.650 ;
        RECT  18.570 1.390 18.690 1.830 ;
        RECT  18.690 1.390 18.930 3.340 ;
        RECT  18.930 2.390 18.940 2.650 ;
        RECT  18.930 2.940 18.970 3.340 ;
        RECT  18.930 1.390 18.970 1.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.720 2.190 2.120 2.630 ;
        RECT  2.120 2.390 2.180 2.630 ;
        RECT  2.180 2.390 2.440 2.650 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  3.500 2.390 3.570 2.650 ;
        RECT  3.570 1.950 3.760 2.650 ;
        RECT  3.760 1.950 3.810 2.640 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.360 5.440 ;
        RECT  0.360 4.480 0.760 5.440 ;
        RECT  0.760 4.640 3.020 5.440 ;
        RECT  3.020 4.480 3.420 5.440 ;
        RECT  3.420 4.640 6.250 5.440 ;
        RECT  6.250 4.480 6.650 5.440 ;
        RECT  6.650 4.640 7.850 5.440 ;
        RECT  7.850 4.480 8.250 5.440 ;
        RECT  11.450 3.410 11.850 3.850 ;
        RECT  11.850 3.610 13.640 3.850 ;
        RECT  13.640 3.410 13.880 3.850 ;
        RECT  13.880 3.410 14.030 3.650 ;
        RECT  14.030 3.280 14.430 3.650 ;
        RECT  8.250 4.640 15.360 5.440 ;
        RECT  14.430 3.410 15.360 3.650 ;
        RECT  15.360 3.410 15.600 5.440 ;
        RECT  15.600 4.640 16.120 5.440 ;
        RECT  16.120 3.390 16.130 5.440 ;
        RECT  16.130 3.270 16.530 5.440 ;
        RECT  16.530 3.390 16.540 5.440 ;
        RECT  16.540 4.640 17.740 5.440 ;
        RECT  17.740 4.480 18.140 5.440 ;
        RECT  18.140 4.640 19.140 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.410 0.400 ;
        RECT  0.410 -0.400 0.830 1.800 ;
        RECT  0.830 1.390 0.900 1.790 ;
        RECT  0.830 -0.400 3.100 0.400 ;
        RECT  3.100 -0.400 3.500 0.560 ;
        RECT  3.500 -0.400 5.870 0.400 ;
        RECT  5.870 -0.400 5.880 0.730 ;
        RECT  5.880 -0.400 6.280 0.850 ;
        RECT  6.280 -0.400 6.290 0.730 ;
        RECT  6.290 -0.400 9.460 0.400 ;
        RECT  9.460 -0.400 9.470 0.730 ;
        RECT  9.470 -0.400 9.870 0.850 ;
        RECT  9.870 -0.400 9.880 0.730 ;
        RECT  9.880 -0.400 11.570 0.400 ;
        RECT  11.570 -0.400 11.580 0.930 ;
        RECT  11.580 -0.400 11.980 1.050 ;
        RECT  11.980 -0.400 11.990 0.930 ;
        RECT  11.990 -0.400 14.270 0.400 ;
        RECT  14.270 -0.400 14.670 0.560 ;
        RECT  14.670 -0.400 17.690 0.400 ;
        RECT  17.690 -0.400 18.090 0.560 ;
        RECT  18.090 -0.400 19.140 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  18.050 0.860 18.290 3.970 ;
        RECT  17.210 0.860 18.050 1.100 ;
        RECT  17.270 3.730 18.050 3.970 ;
        RECT  16.870 3.730 17.270 4.130 ;
        RECT  16.210 2.240 17.250 2.660 ;
        RECT  16.810 0.730 17.210 1.100 ;
        RECT  15.970 1.390 16.210 2.990 ;
        RECT  15.810 1.390 15.970 1.790 ;
        RECT  15.250 2.750 15.970 2.990 ;
        RECT  15.150 2.070 15.550 2.470 ;
        RECT  14.850 2.750 15.250 3.130 ;
        RECT  13.360 2.070 15.150 2.310 ;
        RECT  14.110 2.750 14.850 2.990 ;
        RECT  13.710 2.590 14.110 2.990 ;
        RECT  12.660 0.670 13.540 0.910 ;
        RECT  13.120 1.250 13.360 3.330 ;
        RECT  12.940 1.250 13.120 1.650 ;
        RECT  12.670 3.090 13.120 3.330 ;
        RECT  12.660 2.520 12.840 2.760 ;
        RECT  12.420 0.670 12.660 2.760 ;
        RECT  10.670 1.330 12.420 1.570 ;
        RECT  12.240 2.520 12.420 2.760 ;
        RECT  12.000 2.520 12.240 3.130 ;
        RECT  11.720 1.850 12.120 2.140 ;
        RECT  11.010 2.890 12.000 3.130 ;
        RECT  10.150 1.850 11.720 2.090 ;
        RECT  10.490 2.370 11.400 2.610 ;
        RECT  10.770 2.890 11.010 3.730 ;
        RECT  10.430 0.680 10.670 1.570 ;
        RECT  10.250 2.370 10.490 3.840 ;
        RECT  9.290 3.600 10.250 3.840 ;
        RECT  9.910 1.130 10.150 2.090 ;
        RECT  9.740 2.430 9.970 3.320 ;
        RECT  9.190 1.130 9.910 1.370 ;
        RECT  9.630 2.420 9.740 3.320 ;
        RECT  9.570 1.650 9.630 3.320 ;
        RECT  9.390 1.650 9.570 3.140 ;
        RECT  9.220 1.650 9.390 1.890 ;
        RECT  8.510 2.900 9.390 3.140 ;
        RECT  9.050 3.420 9.290 3.840 ;
        RECT  8.950 0.750 9.190 1.370 ;
        RECT  5.710 3.420 9.050 3.660 ;
        RECT  7.760 0.750 8.950 0.990 ;
        RECT  8.270 2.430 8.510 3.140 ;
        RECT  7.760 1.810 7.990 3.140 ;
        RECT  7.750 0.750 7.760 3.140 ;
        RECT  7.520 0.750 7.750 2.050 ;
        RECT  6.230 2.900 7.750 3.140 ;
        RECT  7.240 2.330 7.470 2.570 ;
        RECT  7.000 1.130 7.240 2.570 ;
        RECT  5.280 1.130 7.000 1.370 ;
        RECT  5.990 2.610 6.230 3.140 ;
        RECT  5.470 2.050 5.710 4.370 ;
        RECT  5.160 2.050 5.470 2.450 ;
        RECT  4.670 4.130 5.470 4.370 ;
        RECT  4.880 0.670 5.280 1.370 ;
        RECT  4.950 2.730 5.190 3.850 ;
        RECT  4.880 2.730 4.950 2.970 ;
        RECT  4.640 1.130 4.880 2.970 ;
        RECT  4.430 3.250 4.670 4.370 ;
        RECT  4.380 3.250 4.430 3.650 ;
        RECT  4.360 3.250 4.380 3.490 ;
        RECT  4.120 1.410 4.360 3.490 ;
        RECT  3.850 0.670 4.250 1.100 ;
        RECT  3.910 3.940 4.150 4.370 ;
        RECT  3.850 1.410 4.120 1.650 ;
        RECT  3.730 3.230 4.120 3.490 ;
        RECT  3.260 3.940 3.910 4.180 ;
        RECT  2.250 0.860 3.850 1.100 ;
        RECT  3.020 3.610 3.260 4.180 ;
        RECT  2.250 3.610 3.020 3.850 ;
        RECT  2.420 4.130 2.500 4.370 ;
        RECT  2.100 4.120 2.420 4.370 ;
        RECT  1.840 0.670 2.250 1.100 ;
        RECT  2.010 3.120 2.250 3.850 ;
        RECT  1.320 4.120 2.100 4.360 ;
        RECT  1.850 3.120 2.010 3.520 ;
        RECT  1.430 0.670 1.510 0.910 ;
        RECT  1.320 0.670 1.430 2.390 ;
        RECT  1.190 0.670 1.320 4.360 ;
        RECT  1.110 0.670 1.190 0.910 ;
        RECT  1.080 2.070 1.190 4.360 ;
    END
END SDFFNSRXL

MACRO SDFFNSRX4
    CLASS CORE ;
    FOREIGN SDFFNSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNSRXL ;
    SIZE 26.400 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.420 3.990 7.820 4.360 ;
        RECT  7.820 4.120 11.300 4.360 ;
        RECT  11.300 3.940 11.760 4.360 ;
        RECT  11.760 3.940 16.290 4.180 ;
        RECT  16.290 3.940 16.820 4.310 ;
        RECT  16.820 3.940 16.970 4.300 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.950 2.850 3.210 ;
        RECT  2.850 2.150 3.090 3.210 ;
        RECT  3.090 2.950 3.100 3.210 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.780 2.500 0.860 2.900 ;
        RECT  0.860 2.390 1.120 2.900 ;
        RECT  1.120 2.500 1.180 2.900 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.350 2.380 9.820 2.810 ;
        RECT  9.820 2.400 9.890 2.800 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  23.210 1.820 23.330 3.220 ;
        RECT  23.330 1.590 23.340 3.220 ;
        RECT  23.340 1.390 23.650 3.220 ;
        RECT  23.650 1.390 23.740 3.150 ;
        RECT  23.740 1.590 23.750 2.950 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  24.530 1.820 24.870 3.220 ;
        RECT  24.870 1.590 24.880 3.220 ;
        RECT  24.880 1.390 24.970 3.220 ;
        RECT  24.970 1.390 25.080 3.160 ;
        RECT  25.080 1.390 25.280 3.150 ;
        RECT  25.280 1.590 25.290 2.820 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.810 2.580 2.110 2.820 ;
        RECT  2.110 2.400 2.180 2.820 ;
        RECT  2.180 2.390 2.350 2.820 ;
        RECT  2.350 2.390 2.440 2.650 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  3.490 1.820 3.850 2.360 ;
        RECT  3.850 1.950 4.030 2.350 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.780 5.440 ;
        RECT  0.780 4.480 1.180 5.440 ;
        RECT  1.180 4.640 3.120 5.440 ;
        RECT  3.120 4.480 3.520 5.440 ;
        RECT  3.520 4.640 6.750 5.440 ;
        RECT  6.750 4.480 7.150 5.440 ;
        RECT  7.150 4.640 12.210 5.440 ;
        RECT  12.210 4.480 12.610 5.440 ;
        RECT  12.610 4.640 14.810 5.440 ;
        RECT  14.810 4.480 15.210 5.440 ;
        RECT  15.210 4.640 17.880 5.440 ;
        RECT  17.880 3.230 17.890 5.440 ;
        RECT  17.890 3.110 18.290 5.440 ;
        RECT  18.290 3.230 18.300 5.440 ;
        RECT  18.300 4.640 19.860 5.440 ;
        RECT  19.860 3.500 19.870 5.440 ;
        RECT  19.870 3.300 20.270 5.440 ;
        RECT  20.270 3.500 20.280 5.440 ;
        RECT  20.280 4.640 22.720 5.440 ;
        RECT  22.720 4.210 22.730 5.440 ;
        RECT  22.730 4.010 23.130 5.440 ;
        RECT  23.130 4.210 23.140 5.440 ;
        RECT  23.140 4.640 24.120 5.440 ;
        RECT  24.120 4.210 24.130 5.440 ;
        RECT  24.130 4.010 24.530 5.440 ;
        RECT  24.530 4.210 24.540 5.440 ;
        RECT  24.540 4.640 25.540 5.440 ;
        RECT  25.540 4.210 25.550 5.440 ;
        RECT  25.550 4.010 25.950 5.440 ;
        RECT  25.950 4.210 25.960 5.440 ;
        RECT  25.960 4.640 26.400 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 0.850 0.730 ;
        RECT  0.850 -0.400 1.250 0.930 ;
        RECT  1.250 -0.400 1.260 0.730 ;
        RECT  1.260 -0.400 3.400 0.400 ;
        RECT  3.400 -0.400 3.800 0.560 ;
        RECT  3.800 -0.400 6.580 0.400 ;
        RECT  6.580 -0.400 6.590 0.730 ;
        RECT  6.590 -0.400 6.990 0.850 ;
        RECT  6.990 -0.400 7.000 0.730 ;
        RECT  7.000 -0.400 10.000 0.400 ;
        RECT  10.000 -0.400 10.010 0.800 ;
        RECT  10.010 -0.400 10.410 0.920 ;
        RECT  10.410 -0.400 10.420 0.800 ;
        RECT  10.420 -0.400 12.080 0.400 ;
        RECT  12.080 -0.400 12.090 0.940 ;
        RECT  12.090 -0.400 12.490 1.060 ;
        RECT  12.490 -0.400 12.500 0.940 ;
        RECT  12.500 -0.400 14.640 0.400 ;
        RECT  14.640 -0.400 14.650 0.820 ;
        RECT  14.650 -0.400 15.050 0.940 ;
        RECT  15.050 -0.400 15.060 0.820 ;
        RECT  15.060 -0.400 17.580 0.400 ;
        RECT  17.580 -0.400 17.590 1.060 ;
        RECT  17.590 -0.400 17.990 1.260 ;
        RECT  17.990 -0.400 18.000 1.060 ;
        RECT  18.000 -0.400 22.720 0.400 ;
        RECT  22.720 -0.400 22.730 0.910 ;
        RECT  22.730 -0.400 23.130 1.110 ;
        RECT  23.130 -0.400 23.140 0.910 ;
        RECT  23.140 -0.400 24.120 0.400 ;
        RECT  24.120 -0.400 24.130 0.910 ;
        RECT  24.130 -0.400 24.530 1.110 ;
        RECT  24.530 -0.400 24.540 0.910 ;
        RECT  24.540 -0.400 25.540 0.400 ;
        RECT  25.540 -0.400 25.550 0.910 ;
        RECT  25.550 -0.400 25.950 1.110 ;
        RECT  25.950 -0.400 25.960 0.910 ;
        RECT  25.960 -0.400 26.400 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  25.560 2.180 25.800 3.730 ;
        RECT  22.940 3.490 25.560 3.730 ;
        RECT  22.700 1.550 22.940 3.730 ;
        RECT  22.230 1.550 22.700 1.790 ;
        RECT  21.860 3.330 22.700 3.730 ;
        RECT  22.020 2.130 22.420 2.530 ;
        RECT  21.990 1.390 22.230 1.790 ;
        RECT  21.670 2.140 22.020 2.530 ;
        RECT  21.390 0.680 21.790 0.960 ;
        RECT  21.490 1.540 21.670 3.020 ;
        RECT  21.430 1.540 21.490 3.930 ;
        RECT  21.030 1.540 21.430 1.780 ;
        RECT  21.090 2.780 21.430 3.930 ;
        RECT  20.270 0.680 21.390 0.920 ;
        RECT  20.910 2.060 21.150 2.500 ;
        RECT  19.050 2.780 21.090 3.020 ;
        RECT  20.630 1.200 21.030 1.780 ;
        RECT  16.600 2.060 20.910 2.300 ;
        RECT  19.510 1.540 20.630 1.780 ;
        RECT  19.870 0.680 20.270 1.260 ;
        RECT  18.750 0.680 19.870 0.920 ;
        RECT  19.110 1.230 19.510 1.780 ;
        RECT  18.890 2.780 19.050 3.920 ;
        RECT  18.650 2.580 18.890 3.920 ;
        RECT  18.590 0.680 18.750 1.490 ;
        RECT  17.530 2.580 18.650 2.820 ;
        RECT  18.510 0.680 18.590 1.780 ;
        RECT  18.350 1.090 18.510 1.780 ;
        RECT  17.150 1.540 18.350 1.780 ;
        RECT  17.370 3.420 17.610 4.360 ;
        RECT  17.290 2.580 17.530 3.140 ;
        RECT  11.180 3.420 17.370 3.660 ;
        RECT  17.130 2.860 17.290 3.140 ;
        RECT  16.910 0.930 17.150 1.780 ;
        RECT  15.430 2.900 17.130 3.140 ;
        RECT  16.360 0.830 16.600 2.300 ;
        RECT  15.990 0.830 16.360 1.070 ;
        RECT  16.110 1.920 16.360 2.300 ;
        RECT  15.710 1.920 16.110 2.620 ;
        RECT  15.640 1.400 16.070 1.640 ;
        RECT  14.210 1.920 15.710 2.160 ;
        RECT  15.400 1.230 15.640 1.640 ;
        RECT  15.190 2.440 15.430 3.140 ;
        RECT  14.370 1.230 15.400 1.470 ;
        RECT  15.030 2.440 15.190 2.680 ;
        RECT  14.130 0.670 14.370 1.470 ;
        RECT  13.970 1.750 14.210 3.140 ;
        RECT  13.170 0.670 14.130 0.910 ;
        RECT  13.690 1.750 13.970 1.990 ;
        RECT  13.480 2.900 13.970 3.140 ;
        RECT  13.450 1.190 13.690 1.990 ;
        RECT  13.170 2.270 13.640 2.510 ;
        RECT  12.930 0.670 13.170 2.910 ;
        RECT  11.590 1.340 12.930 1.580 ;
        RECT  11.860 2.670 12.930 2.910 ;
        RECT  10.970 1.860 12.650 2.100 ;
        RECT  11.540 2.670 11.860 3.140 ;
        RECT  11.350 0.680 11.590 1.580 ;
        RECT  11.460 2.900 11.540 3.140 ;
        RECT  10.910 0.680 11.350 0.920 ;
        RECT  10.940 3.080 11.180 3.660 ;
        RECT  10.730 1.200 10.970 2.100 ;
        RECT  10.450 3.080 10.940 3.320 ;
        RECT  9.770 1.200 10.730 1.440 ;
        RECT  8.340 3.600 10.660 3.840 ;
        RECT  10.210 1.720 10.450 3.320 ;
        RECT  10.050 1.720 10.210 1.960 ;
        RECT  9.030 3.080 10.210 3.320 ;
        RECT  9.530 1.200 9.770 1.990 ;
        RECT  8.570 1.750 9.530 1.990 ;
        RECT  9.010 0.670 9.250 1.470 ;
        RECT  8.790 2.370 9.030 3.320 ;
        RECT  7.730 0.670 9.010 0.910 ;
        RECT  8.510 1.190 8.570 1.990 ;
        RECT  8.270 1.190 8.510 3.100 ;
        RECT  8.100 3.470 8.340 3.840 ;
        RECT  8.170 1.190 8.270 1.430 ;
        RECT  8.090 2.860 8.270 3.100 ;
        RECT  6.310 3.470 8.100 3.710 ;
        RECT  7.690 2.860 8.090 3.190 ;
        RECT  7.750 1.710 7.990 2.140 ;
        RECT  7.110 1.710 7.750 1.950 ;
        RECT  7.490 0.670 7.730 1.360 ;
        RECT  6.830 2.860 7.690 3.100 ;
        RECT  6.870 1.190 7.110 1.950 ;
        RECT  5.870 1.190 6.870 1.430 ;
        RECT  6.590 2.300 6.830 3.100 ;
        RECT  6.070 1.820 6.310 4.370 ;
        RECT  5.680 1.820 6.070 2.060 ;
        RECT  5.270 4.130 6.070 4.370 ;
        RECT  5.470 0.670 5.870 1.430 ;
        RECT  5.550 2.530 5.790 3.850 ;
        RECT  5.400 2.530 5.550 2.770 ;
        RECT  5.400 1.190 5.470 1.430 ;
        RECT  5.160 1.190 5.400 2.770 ;
        RECT  5.080 3.080 5.270 4.370 ;
        RECT  4.870 0.670 5.110 0.910 ;
        RECT  5.030 3.070 5.080 4.370 ;
        RECT  4.640 3.070 5.030 3.460 ;
        RECT  4.630 0.670 4.870 1.100 ;
        RECT  4.510 3.730 4.750 4.130 ;
        RECT  4.480 1.410 4.640 3.460 ;
        RECT  2.630 0.860 4.630 1.100 ;
        RECT  3.590 3.730 4.510 3.970 ;
        RECT  4.400 1.410 4.480 3.450 ;
        RECT  4.220 1.410 4.400 1.650 ;
        RECT  3.930 2.990 4.400 3.450 ;
        RECT  3.350 3.600 3.590 3.970 ;
        RECT  2.450 3.600 3.350 3.840 ;
        RECT  1.690 4.120 2.780 4.360 ;
        RECT  2.390 0.860 2.630 1.650 ;
        RECT  2.210 3.100 2.450 3.840 ;
        RECT  2.230 1.250 2.390 1.650 ;
        RECT  2.050 3.100 2.210 3.500 ;
        RECT  1.450 3.180 1.690 4.360 ;
        RECT  0.570 1.860 1.590 2.100 ;
        RECT  0.410 3.180 1.450 3.420 ;
        RECT  0.410 1.370 0.570 2.100 ;
        RECT  0.170 1.370 0.410 3.420 ;
    END
END SDFFNSRX4

MACRO SDFFNSRX2
    CLASS CORE ;
    FOREIGN SDFFNSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNSRXL ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.520 3.940 6.920 4.370 ;
        RECT  6.920 3.940 7.950 4.180 ;
        RECT  7.950 3.940 8.190 4.360 ;
        RECT  8.190 4.120 10.400 4.360 ;
        RECT  10.400 4.120 10.770 4.370 ;
        RECT  10.770 4.130 13.990 4.370 ;
        RECT  13.990 4.030 14.390 4.370 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.430 2.280 2.580 2.680 ;
        RECT  2.580 2.280 2.820 3.190 ;
        RECT  2.820 2.280 2.830 2.680 ;
        RECT  2.820 2.950 2.840 3.190 ;
        RECT  2.840 2.950 3.100 3.210 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.680 0.860 3.200 ;
        RECT  0.860 2.680 0.920 3.210 ;
        RECT  0.920 2.950 1.120 3.210 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.120 1.770 8.770 2.190 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.360 2.640 17.520 3.210 ;
        RECT  17.520 1.160 17.760 3.210 ;
        RECT  17.760 1.160 18.110 1.560 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.680 2.950 18.790 3.210 ;
        RECT  18.790 2.940 19.130 3.220 ;
        RECT  19.130 2.940 19.390 4.160 ;
        RECT  19.230 0.950 19.390 1.350 ;
        RECT  19.390 0.950 19.530 4.160 ;
        RECT  19.530 0.950 19.630 4.150 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.330 2.270 1.910 2.670 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  3.230 1.950 3.470 2.630 ;
        RECT  3.470 2.390 3.500 2.630 ;
        RECT  3.500 2.390 3.760 2.650 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 2.750 5.440 ;
        RECT  2.750 4.480 3.150 5.440 ;
        RECT  3.150 4.640 5.840 5.440 ;
        RECT  5.840 4.480 6.240 5.440 ;
        RECT  6.240 4.640 7.270 5.440 ;
        RECT  7.270 4.480 7.670 5.440 ;
        RECT  11.080 3.510 11.480 3.850 ;
        RECT  11.480 3.610 13.290 3.850 ;
        RECT  13.290 3.470 13.530 3.850 ;
        RECT  7.670 4.640 14.690 5.440 ;
        RECT  13.530 3.470 14.690 3.710 ;
        RECT  14.690 3.470 14.930 5.440 ;
        RECT  14.930 4.640 15.810 5.440 ;
        RECT  15.810 3.730 15.820 5.440 ;
        RECT  15.820 3.530 16.220 5.440 ;
        RECT  16.220 3.730 16.230 5.440 ;
        RECT  16.230 4.640 18.300 5.440 ;
        RECT  18.300 4.360 18.310 5.440 ;
        RECT  18.310 4.160 18.710 5.440 ;
        RECT  18.710 4.360 18.720 5.440 ;
        RECT  18.720 4.640 19.800 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.440 0.400 ;
        RECT  0.440 -0.400 0.450 0.750 ;
        RECT  0.450 -0.400 0.850 0.870 ;
        RECT  0.850 -0.400 0.860 0.750 ;
        RECT  0.860 -0.400 2.750 0.400 ;
        RECT  2.750 -0.400 3.150 0.560 ;
        RECT  3.150 -0.400 5.870 0.400 ;
        RECT  5.870 -0.400 5.880 0.730 ;
        RECT  5.880 -0.400 6.280 0.850 ;
        RECT  6.280 -0.400 6.290 0.730 ;
        RECT  6.290 -0.400 8.920 0.400 ;
        RECT  8.920 -0.400 8.930 0.730 ;
        RECT  8.930 -0.400 9.330 0.850 ;
        RECT  9.330 -0.400 9.340 0.730 ;
        RECT  9.340 -0.400 11.170 0.400 ;
        RECT  11.170 -0.400 11.180 0.750 ;
        RECT  11.180 -0.400 11.580 0.870 ;
        RECT  11.580 -0.400 11.590 0.750 ;
        RECT  11.590 -0.400 13.750 0.400 ;
        RECT  13.750 -0.400 14.150 0.560 ;
        RECT  14.150 -0.400 16.910 0.400 ;
        RECT  16.910 -0.400 17.310 0.560 ;
        RECT  17.310 -0.400 18.460 0.400 ;
        RECT  18.460 -0.400 18.470 1.220 ;
        RECT  18.470 -0.400 18.870 1.710 ;
        RECT  18.870 -0.400 18.880 1.220 ;
        RECT  18.880 -0.400 19.800 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  18.690 2.240 19.090 2.640 ;
        RECT  18.320 2.400 18.690 2.640 ;
        RECT  18.080 2.400 18.320 3.730 ;
        RECT  17.050 3.490 18.080 3.730 ;
        RECT  17.000 1.300 17.240 1.700 ;
        RECT  17.000 3.490 17.050 3.890 ;
        RECT  16.760 1.300 17.000 3.890 ;
        RECT  16.650 3.490 16.760 3.890 ;
        RECT  16.400 0.750 16.480 1.150 ;
        RECT  15.720 2.270 16.480 2.670 ;
        RECT  16.080 0.740 16.400 1.150 ;
        RECT  14.960 0.740 16.080 0.980 ;
        RECT  15.480 1.280 15.720 3.170 ;
        RECT  15.320 1.280 15.480 1.520 ;
        RECT  13.790 2.930 15.480 3.170 ;
        RECT  14.800 1.790 15.200 2.190 ;
        RECT  14.640 0.740 14.960 1.150 ;
        RECT  13.040 1.850 14.800 2.090 ;
        RECT  14.560 0.750 14.640 1.150 ;
        RECT  13.550 2.610 13.790 3.170 ;
        RECT  13.380 2.610 13.550 2.850 ;
        RECT  12.260 0.730 13.320 0.970 ;
        RECT  13.000 1.330 13.040 2.090 ;
        RECT  12.760 1.330 13.000 3.330 ;
        RECT  12.620 1.330 12.760 1.570 ;
        RECT  12.380 3.090 12.760 3.330 ;
        RECT  12.260 2.520 12.480 2.760 ;
        RECT  12.020 0.730 12.260 2.760 ;
        RECT  10.640 1.150 12.020 1.390 ;
        RECT  11.910 2.520 12.020 2.760 ;
        RECT  11.670 2.520 11.910 3.130 ;
        RECT  11.320 1.850 11.720 2.140 ;
        RECT  10.640 2.890 11.670 3.130 ;
        RECT  9.960 1.850 11.320 2.090 ;
        RECT  10.010 2.370 11.000 2.610 ;
        RECT  10.480 1.150 10.640 1.570 ;
        RECT  10.400 2.890 10.640 3.830 ;
        RECT  10.240 0.670 10.480 1.570 ;
        RECT  9.770 2.370 10.010 3.840 ;
        RECT  9.720 1.130 9.960 2.090 ;
        RECT  8.710 3.600 9.770 3.840 ;
        RECT  8.550 1.130 9.720 1.370 ;
        RECT  9.440 2.430 9.480 3.320 ;
        RECT  9.200 1.650 9.440 3.320 ;
        RECT  9.040 1.650 9.200 1.890 ;
        RECT  8.990 2.900 9.200 3.320 ;
        RECT  8.260 2.900 8.990 3.140 ;
        RECT  8.470 3.420 8.710 3.840 ;
        RECT  8.310 1.130 8.550 1.430 ;
        RECT  5.540 3.420 8.470 3.660 ;
        RECT  7.740 1.190 8.310 1.430 ;
        RECT  8.020 2.510 8.260 3.140 ;
        RECT  7.500 1.190 7.740 3.140 ;
        RECT  7.420 1.190 7.500 1.430 ;
        RECT  6.060 2.900 7.500 3.140 ;
        RECT  6.980 1.740 7.220 2.190 ;
        RECT  6.080 1.740 6.980 1.980 ;
        RECT  5.840 1.130 6.080 1.980 ;
        RECT  5.820 2.490 6.060 3.140 ;
        RECT  4.940 1.130 5.840 1.370 ;
        RECT  5.300 1.740 5.540 4.370 ;
        RECT  5.160 1.740 5.300 2.140 ;
        RECT  4.460 4.130 5.300 4.370 ;
        RECT  4.980 3.450 5.020 3.850 ;
        RECT  4.880 2.730 4.980 3.850 ;
        RECT  4.880 0.740 4.940 1.370 ;
        RECT  4.740 0.740 4.880 3.850 ;
        RECT  4.640 0.740 4.740 2.970 ;
        RECT  4.540 0.740 4.640 1.140 ;
        RECT  4.370 3.250 4.460 4.370 ;
        RECT  4.220 1.410 4.370 4.370 ;
        RECT  4.130 1.410 4.220 3.650 ;
        RECT  3.630 1.410 4.130 1.650 ;
        RECT  3.560 3.250 4.130 3.650 ;
        RECT  3.630 0.670 4.030 1.100 ;
        RECT  3.700 3.940 3.940 4.370 ;
        RECT  3.260 3.940 3.700 4.180 ;
        RECT  2.260 0.860 3.630 1.100 ;
        RECT  3.020 3.610 3.260 4.180 ;
        RECT  2.020 3.610 3.020 3.850 ;
        RECT  2.020 0.860 2.260 1.750 ;
        RECT  1.090 4.130 2.180 4.370 ;
        RECT  1.710 1.350 2.020 1.750 ;
        RECT  1.780 3.340 2.020 3.850 ;
        RECT  1.620 3.340 1.780 3.580 ;
        RECT  1.370 0.670 1.730 0.910 ;
        RECT  1.130 0.670 1.370 1.390 ;
        RECT  0.930 1.150 1.130 1.390 ;
        RECT  0.850 3.940 1.090 4.370 ;
        RECT  0.690 1.150 0.930 2.360 ;
        RECT  0.400 3.940 0.850 4.180 ;
        RECT  0.400 2.120 0.690 2.360 ;
        RECT  0.160 2.120 0.400 4.180 ;
    END
END SDFFNSRX2

MACRO SDFFNSRX1
    CLASS CORE ;
    FOREIGN SDFFNSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNSRXL ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.520 4.130 6.650 4.370 ;
        RECT  6.650 3.940 6.920 4.370 ;
        RECT  6.920 3.940 7.950 4.180 ;
        RECT  7.950 3.940 8.190 4.360 ;
        RECT  8.190 4.120 10.400 4.360 ;
        RECT  10.400 4.120 10.770 4.370 ;
        RECT  10.770 4.130 13.990 4.370 ;
        RECT  13.990 4.030 14.390 4.370 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.420 2.280 2.580 2.680 ;
        RECT  2.580 2.280 2.820 3.190 ;
        RECT  2.820 2.950 2.840 3.190 ;
        RECT  2.840 2.950 3.100 3.210 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.680 0.860 3.200 ;
        RECT  0.860 2.680 0.920 3.210 ;
        RECT  0.920 2.950 1.120 3.210 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.120 1.770 8.670 2.190 ;
        RECT  8.670 1.780 8.760 2.180 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.160 0.740 16.400 3.090 ;
        RECT  16.400 0.740 16.700 0.980 ;
        RECT  16.700 0.710 16.950 0.980 ;
        RECT  16.950 0.710 16.960 0.970 ;
        RECT  16.400 2.850 17.100 3.090 ;
        RECT  16.960 0.730 17.140 0.970 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.570 2.970 18.690 3.370 ;
        RECT  18.680 2.390 18.690 2.650 ;
        RECT  18.570 1.320 18.690 1.830 ;
        RECT  18.690 1.320 18.930 3.370 ;
        RECT  18.930 2.390 18.940 2.650 ;
        RECT  18.930 2.970 18.970 3.370 ;
        RECT  18.930 1.320 18.970 1.960 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.320 2.250 1.330 2.660 ;
        RECT  1.330 2.040 1.770 2.660 ;
        RECT  1.770 2.250 1.780 2.660 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  3.230 1.950 3.470 2.630 ;
        RECT  3.470 2.390 3.500 2.630 ;
        RECT  3.500 2.390 3.760 2.650 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 2.750 5.440 ;
        RECT  2.750 4.480 3.150 5.440 ;
        RECT  3.150 4.640 5.840 5.440 ;
        RECT  5.840 4.480 6.240 5.440 ;
        RECT  6.240 4.640 7.270 5.440 ;
        RECT  7.270 4.480 7.670 5.440 ;
        RECT  11.080 3.520 11.480 3.850 ;
        RECT  11.480 3.610 13.290 3.850 ;
        RECT  13.290 3.470 13.530 3.850 ;
        RECT  7.670 4.640 14.690 5.440 ;
        RECT  13.530 3.470 14.690 3.710 ;
        RECT  14.690 3.470 14.930 5.440 ;
        RECT  14.930 4.640 15.870 5.440 ;
        RECT  15.870 4.050 15.880 5.440 ;
        RECT  15.880 3.930 16.280 5.440 ;
        RECT  16.280 4.050 16.290 5.440 ;
        RECT  16.290 4.640 17.530 5.440 ;
        RECT  17.530 4.480 17.930 5.440 ;
        RECT  17.930 4.640 19.140 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.440 0.400 ;
        RECT  0.440 -0.400 0.450 0.750 ;
        RECT  0.450 -0.400 0.850 0.870 ;
        RECT  0.850 -0.400 0.860 0.750 ;
        RECT  0.860 -0.400 2.890 0.400 ;
        RECT  2.890 -0.400 3.290 0.560 ;
        RECT  3.290 -0.400 5.870 0.400 ;
        RECT  5.870 -0.400 5.880 0.730 ;
        RECT  5.880 -0.400 6.280 0.850 ;
        RECT  6.280 -0.400 6.290 0.730 ;
        RECT  6.290 -0.400 8.920 0.400 ;
        RECT  8.920 -0.400 8.930 0.730 ;
        RECT  8.930 -0.400 9.330 0.850 ;
        RECT  9.330 -0.400 9.340 0.730 ;
        RECT  9.340 -0.400 11.170 0.400 ;
        RECT  11.170 -0.400 11.180 0.930 ;
        RECT  11.180 -0.400 11.580 1.050 ;
        RECT  11.580 -0.400 11.590 0.930 ;
        RECT  11.590 -0.400 13.740 0.400 ;
        RECT  13.740 -0.400 14.140 0.560 ;
        RECT  14.140 -0.400 17.630 0.400 ;
        RECT  17.630 -0.400 17.640 1.070 ;
        RECT  17.640 -0.400 18.040 1.270 ;
        RECT  18.040 -0.400 18.050 1.070 ;
        RECT  18.050 -0.400 19.140 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  18.180 2.180 18.320 2.580 ;
        RECT  18.160 2.180 18.180 4.170 ;
        RECT  17.940 1.550 18.160 4.170 ;
        RECT  17.920 1.550 17.940 2.580 ;
        RECT  17.040 3.930 17.940 4.170 ;
        RECT  17.080 1.550 17.920 1.790 ;
        RECT  17.380 2.170 17.620 3.610 ;
        RECT  17.280 2.170 17.380 2.570 ;
        RECT  15.780 3.370 17.380 3.610 ;
        RECT  16.680 1.390 17.080 1.790 ;
        RECT  16.640 3.930 17.040 4.330 ;
        RECT  15.540 1.490 15.780 3.610 ;
        RECT  15.520 1.490 15.540 1.730 ;
        RECT  13.820 2.930 15.540 3.170 ;
        RECT  15.120 1.330 15.520 1.730 ;
        RECT  14.840 2.160 15.240 2.560 ;
        RECT  13.040 2.160 14.840 2.400 ;
        RECT  13.580 2.680 13.820 3.170 ;
        RECT  13.420 2.680 13.580 2.920 ;
        RECT  12.240 0.730 13.220 0.970 ;
        RECT  13.000 1.300 13.040 2.400 ;
        RECT  12.760 1.300 13.000 3.330 ;
        RECT  12.520 1.300 12.760 1.540 ;
        RECT  12.380 3.090 12.760 3.330 ;
        RECT  12.240 2.520 12.480 2.760 ;
        RECT  12.000 0.730 12.240 2.760 ;
        RECT  11.900 0.730 12.000 1.570 ;
        RECT  11.910 2.520 12.000 2.760 ;
        RECT  11.670 2.520 11.910 3.130 ;
        RECT  10.480 1.330 11.900 1.570 ;
        RECT  11.320 1.850 11.720 2.110 ;
        RECT  10.640 2.890 11.670 3.130 ;
        RECT  9.960 1.850 11.320 2.090 ;
        RECT  10.010 2.370 11.000 2.610 ;
        RECT  10.400 2.890 10.640 3.830 ;
        RECT  10.240 0.680 10.480 1.570 ;
        RECT  9.770 2.370 10.010 3.840 ;
        RECT  9.720 1.130 9.960 2.090 ;
        RECT  8.710 3.600 9.770 3.840 ;
        RECT  8.550 1.130 9.720 1.370 ;
        RECT  9.440 2.430 9.480 3.320 ;
        RECT  9.200 1.650 9.440 3.320 ;
        RECT  9.030 1.650 9.200 1.890 ;
        RECT  8.990 2.900 9.200 3.320 ;
        RECT  8.260 2.900 8.990 3.140 ;
        RECT  8.470 3.420 8.710 3.840 ;
        RECT  8.310 1.130 8.550 1.410 ;
        RECT  5.540 3.420 8.470 3.660 ;
        RECT  7.740 1.170 8.310 1.410 ;
        RECT  8.020 2.510 8.260 3.140 ;
        RECT  7.500 1.170 7.740 3.140 ;
        RECT  7.420 1.170 7.500 1.410 ;
        RECT  6.060 2.900 7.500 3.140 ;
        RECT  6.980 1.740 7.220 2.190 ;
        RECT  6.080 1.740 6.980 1.980 ;
        RECT  5.840 1.130 6.080 1.980 ;
        RECT  5.820 2.610 6.060 3.140 ;
        RECT  4.940 1.130 5.840 1.370 ;
        RECT  5.300 1.740 5.540 4.360 ;
        RECT  5.160 1.740 5.300 2.140 ;
        RECT  4.460 4.120 5.300 4.360 ;
        RECT  4.980 3.440 5.020 3.840 ;
        RECT  4.880 2.730 4.980 3.840 ;
        RECT  4.880 0.740 4.940 1.370 ;
        RECT  4.740 0.740 4.880 3.840 ;
        RECT  4.640 0.740 4.740 2.970 ;
        RECT  4.540 0.740 4.640 1.140 ;
        RECT  4.370 3.250 4.460 4.360 ;
        RECT  4.220 1.410 4.370 4.360 ;
        RECT  4.130 1.410 4.220 3.650 ;
        RECT  3.630 1.410 4.130 1.650 ;
        RECT  3.560 3.250 4.130 3.650 ;
        RECT  3.880 0.670 4.030 0.910 ;
        RECT  3.700 3.940 3.940 4.370 ;
        RECT  3.630 0.670 3.880 1.100 ;
        RECT  3.260 3.940 3.700 4.180 ;
        RECT  2.260 0.860 3.630 1.100 ;
        RECT  3.020 3.610 3.260 4.180 ;
        RECT  2.020 3.610 3.020 3.850 ;
        RECT  1.090 4.130 2.320 4.370 ;
        RECT  2.020 0.860 2.260 1.590 ;
        RECT  1.950 1.350 2.020 1.590 ;
        RECT  1.780 3.340 2.020 3.850 ;
        RECT  1.710 1.350 1.950 1.750 ;
        RECT  1.620 3.340 1.780 3.580 ;
        RECT  1.370 0.670 1.730 0.910 ;
        RECT  1.130 0.670 1.370 1.390 ;
        RECT  0.930 1.150 1.130 1.390 ;
        RECT  0.850 3.940 1.090 4.370 ;
        RECT  0.690 1.150 0.930 2.360 ;
        RECT  0.400 3.940 0.850 4.180 ;
        RECT  0.400 2.120 0.690 2.360 ;
        RECT  0.160 2.120 0.400 4.180 ;
    END
END SDFFNSRX1

MACRO SDFFNSXL
    CLASS CORE ;
    FOREIGN SDFFNSXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  12.740 4.070 12.750 4.330 ;
        RECT  12.750 4.060 13.000 4.330 ;
        RECT  13.000 4.060 13.100 4.300 ;
        RECT  13.100 3.740 13.340 4.300 ;
        RECT  13.340 3.740 13.500 4.140 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.380 2.080 3.390 2.650 ;
        RECT  3.390 2.020 3.790 2.650 ;
        RECT  3.790 2.080 3.800 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.470 1.700 1.870 2.300 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.470 3.520 14.720 3.950 ;
        RECT  14.720 3.510 14.870 3.950 ;
        RECT  14.530 0.690 14.930 1.100 ;
        RECT  14.870 3.510 14.980 3.770 ;
        RECT  14.930 0.860 15.290 1.100 ;
        RECT  14.980 3.520 15.430 3.760 ;
        RECT  15.290 0.860 15.430 1.280 ;
        RECT  15.430 0.860 15.670 3.760 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.000 1.280 16.300 3.570 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.130 1.690 4.680 2.090 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.290 0.800 2.690 ;
        RECT  0.800 2.280 1.130 2.700 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.270 5.440 ;
        RECT  0.270 4.480 0.670 5.440 ;
        RECT  0.670 4.640 3.460 5.440 ;
        RECT  3.460 4.270 3.470 5.440 ;
        RECT  3.470 4.150 3.870 5.440 ;
        RECT  3.870 4.270 3.880 5.440 ;
        RECT  3.880 4.640 6.700 5.440 ;
        RECT  6.700 4.480 7.100 5.440 ;
        RECT  7.100 4.640 8.220 5.440 ;
        RECT  8.220 4.310 8.230 5.440 ;
        RECT  8.230 4.190 8.630 5.440 ;
        RECT  8.630 4.310 8.640 5.440 ;
        RECT  8.640 4.640 9.540 5.440 ;
        RECT  9.540 4.040 9.550 5.440 ;
        RECT  9.550 3.840 9.950 5.440 ;
        RECT  9.950 4.040 9.960 5.440 ;
        RECT  9.960 4.640 11.940 5.440 ;
        RECT  11.940 4.210 11.950 5.440 ;
        RECT  11.950 4.010 12.350 5.440 ;
        RECT  12.350 4.210 12.360 5.440 ;
        RECT  12.360 4.640 13.790 5.440 ;
        RECT  13.790 3.730 14.030 5.440 ;
        RECT  14.030 4.640 15.260 5.440 ;
        RECT  15.260 4.480 15.660 5.440 ;
        RECT  15.660 4.640 16.500 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.020 0.400 ;
        RECT  1.020 -0.400 1.420 0.560 ;
        RECT  1.420 -0.400 3.090 0.400 ;
        RECT  3.090 -0.400 3.490 0.560 ;
        RECT  3.490 -0.400 6.640 0.400 ;
        RECT  6.640 -0.400 6.650 0.750 ;
        RECT  6.650 -0.400 7.050 0.870 ;
        RECT  7.050 -0.400 7.060 0.750 ;
        RECT  7.060 -0.400 9.300 0.400 ;
        RECT  9.300 -0.400 9.310 0.750 ;
        RECT  9.310 -0.400 9.710 0.870 ;
        RECT  9.710 -0.400 9.720 0.750 ;
        RECT  9.720 -0.400 11.570 0.400 ;
        RECT  11.570 -0.400 11.970 0.560 ;
        RECT  11.970 -0.400 13.640 0.400 ;
        RECT  13.640 -0.400 13.650 0.850 ;
        RECT  13.650 -0.400 14.050 1.050 ;
        RECT  14.050 -0.400 14.060 0.850 ;
        RECT  14.060 -0.400 15.260 0.400 ;
        RECT  15.260 -0.400 15.660 0.560 ;
        RECT  15.660 -0.400 16.500 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.940 1.960 15.150 2.370 ;
        RECT  14.930 1.500 14.940 2.370 ;
        RECT  14.690 1.380 14.930 3.210 ;
        RECT  14.680 1.380 14.690 2.110 ;
        RECT  14.530 2.810 14.690 3.210 ;
        RECT  14.530 1.380 14.680 1.780 ;
        RECT  14.090 2.020 14.250 2.420 ;
        RECT  13.850 1.570 14.090 3.210 ;
        RECT  12.710 1.570 13.850 1.810 ;
        RECT  13.230 2.970 13.850 3.210 ;
        RECT  12.830 2.970 13.230 3.370 ;
        RECT  12.530 2.290 12.930 2.690 ;
        RECT  12.310 1.220 12.710 1.810 ;
        RECT  11.510 2.370 12.530 2.610 ;
        RECT  12.030 1.570 12.310 1.810 ;
        RECT  11.790 1.570 12.030 1.970 ;
        RECT  11.270 1.610 11.510 3.760 ;
        RECT  10.770 1.610 11.270 1.850 ;
        RECT  10.830 3.360 11.270 3.760 ;
        RECT  10.250 0.670 11.150 0.910 ;
        RECT  10.250 2.810 10.990 3.050 ;
        RECT  10.530 1.450 10.770 1.850 ;
        RECT  10.010 0.670 10.250 3.050 ;
        RECT  8.870 1.240 10.010 1.480 ;
        RECT  9.570 2.810 10.010 3.050 ;
        RECT  9.490 2.020 9.730 2.420 ;
        RECT  9.330 2.810 9.570 3.390 ;
        RECT  8.820 2.100 9.490 2.340 ;
        RECT  9.110 3.150 9.330 3.390 ;
        RECT  8.910 3.670 9.150 4.070 ;
        RECT  6.350 3.670 8.910 3.910 ;
        RECT  8.630 0.670 8.870 1.480 ;
        RECT  8.580 1.760 8.820 3.400 ;
        RECT  7.860 0.670 8.630 0.910 ;
        RECT  8.350 1.760 8.580 2.000 ;
        RECT  6.870 3.160 8.580 3.400 ;
        RECT  8.110 1.430 8.350 2.000 ;
        RECT  7.950 2.370 8.190 2.770 ;
        RECT  7.580 2.370 7.950 2.610 ;
        RECT  7.340 1.150 7.580 2.610 ;
        RECT  5.710 1.150 7.340 1.390 ;
        RECT  6.630 2.530 6.870 3.400 ;
        RECT  6.110 1.830 6.350 4.140 ;
        RECT  5.950 1.830 6.110 2.070 ;
        RECT  4.510 3.900 6.110 4.140 ;
        RECT  5.710 1.670 5.950 2.070 ;
        RECT  5.590 2.520 5.830 3.500 ;
        RECT  5.430 0.760 5.710 1.390 ;
        RECT  5.430 2.520 5.590 2.760 ;
        RECT  5.310 0.760 5.430 2.760 ;
        RECT  5.190 1.150 5.310 2.760 ;
        RECT  4.830 3.100 5.070 3.500 ;
        RECT  4.430 0.750 4.830 1.150 ;
        RECT  2.670 3.110 4.830 3.350 ;
        RECT  4.270 3.630 4.510 4.140 ;
        RECT  2.570 0.860 4.430 1.100 ;
        RECT  3.190 3.630 4.270 3.870 ;
        RECT  2.890 1.380 3.790 1.620 ;
        RECT  2.950 3.630 3.190 4.370 ;
        RECT  2.890 2.540 2.970 2.830 ;
        RECT  1.850 4.130 2.950 4.370 ;
        RECT  2.650 1.380 2.890 2.830 ;
        RECT  2.430 3.110 2.670 3.850 ;
        RECT  2.260 1.420 2.650 1.830 ;
        RECT  2.570 2.540 2.650 2.830 ;
        RECT  2.330 0.670 2.570 1.100 ;
        RECT  2.110 2.590 2.570 2.830 ;
        RECT  2.270 3.610 2.430 3.850 ;
        RECT  1.750 0.670 2.330 0.910 ;
        RECT  2.140 1.430 2.260 1.830 ;
        RECT  1.870 2.590 2.110 3.110 ;
        RECT  1.710 2.870 1.870 3.110 ;
        RECT  1.610 3.910 1.850 4.370 ;
        RECT  0.570 3.910 1.610 4.150 ;
        RECT  0.400 1.270 0.570 1.670 ;
        RECT  0.400 3.100 0.570 4.150 ;
        RECT  0.330 1.270 0.400 4.150 ;
        RECT  0.160 1.270 0.330 3.690 ;
    END
END SDFFNSXL

MACRO SDFFNSX4
    CLASS CORE ;
    FOREIGN SDFFNSX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNSXL ;
    SIZE 21.780 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.370 4.060 7.990 4.380 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.410 2.010 3.850 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 1.700 1.870 2.260 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.920 1.150 18.930 1.680 ;
        RECT  19.050 2.800 19.250 3.200 ;
        RECT  18.930 0.660 19.250 1.680 ;
        RECT  19.250 0.660 19.330 3.210 ;
        RECT  19.330 1.150 19.340 3.210 ;
        RECT  19.340 1.260 19.670 3.210 ;
        RECT  19.670 1.260 19.690 2.660 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  20.450 0.860 20.470 1.260 ;
        RECT  20.560 2.800 20.570 3.200 ;
        RECT  20.470 0.850 20.570 1.260 ;
        RECT  20.570 0.850 20.930 3.220 ;
        RECT  20.930 1.820 21.010 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.380 1.680 4.530 2.080 ;
        RECT  4.530 1.680 4.780 2.090 ;
        RECT  4.780 1.820 5.080 2.090 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.760 2.170 1.170 2.660 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.280 5.440 ;
        RECT  0.280 4.480 0.680 5.440 ;
        RECT  0.680 4.640 3.510 5.440 ;
        RECT  3.510 4.310 3.520 5.440 ;
        RECT  3.520 4.190 3.920 5.440 ;
        RECT  3.920 4.310 3.930 5.440 ;
        RECT  3.930 4.640 6.860 5.440 ;
        RECT  6.860 4.170 7.100 5.440 ;
        RECT  7.100 4.640 8.310 5.440 ;
        RECT  8.310 4.310 8.320 5.440 ;
        RECT  8.320 4.190 8.720 5.440 ;
        RECT  8.720 4.310 8.730 5.440 ;
        RECT  8.730 4.640 9.650 5.440 ;
        RECT  9.650 4.030 9.660 5.440 ;
        RECT  9.660 3.830 10.060 5.440 ;
        RECT  10.060 4.030 10.070 5.440 ;
        RECT  10.070 4.640 12.190 5.440 ;
        RECT  12.190 3.630 12.590 5.440 ;
        RECT  12.590 4.640 14.040 5.440 ;
        RECT  14.040 4.010 14.440 5.440 ;
        RECT  14.440 4.640 15.550 5.440 ;
        RECT  15.550 3.490 15.950 5.440 ;
        RECT  15.950 4.640 16.980 5.440 ;
        RECT  16.980 3.690 16.990 5.440 ;
        RECT  16.990 3.490 17.390 5.440 ;
        RECT  17.390 3.690 17.400 5.440 ;
        RECT  17.400 4.640 18.430 5.440 ;
        RECT  18.430 4.010 18.830 5.440 ;
        RECT  18.830 4.640 19.810 5.440 ;
        RECT  19.810 4.210 19.820 5.440 ;
        RECT  19.820 4.010 20.220 5.440 ;
        RECT  20.220 4.210 20.230 5.440 ;
        RECT  20.230 4.640 21.200 5.440 ;
        RECT  21.200 4.210 21.210 5.440 ;
        RECT  21.210 4.010 21.610 5.440 ;
        RECT  21.610 4.210 21.620 5.440 ;
        RECT  21.620 4.640 21.780 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.180 0.400 ;
        RECT  1.180 -0.400 1.580 0.560 ;
        RECT  1.580 -0.400 3.340 0.400 ;
        RECT  3.340 -0.400 3.740 0.560 ;
        RECT  3.740 -0.400 6.890 0.400 ;
        RECT  6.890 -0.400 6.900 1.000 ;
        RECT  6.900 -0.400 7.300 1.120 ;
        RECT  7.300 -0.400 7.310 1.000 ;
        RECT  7.310 -0.400 9.790 0.400 ;
        RECT  9.790 -0.400 9.800 0.910 ;
        RECT  9.800 -0.400 10.200 1.110 ;
        RECT  10.200 -0.400 10.210 0.910 ;
        RECT  10.210 -0.400 12.420 0.400 ;
        RECT  12.420 -0.400 12.820 0.560 ;
        RECT  12.820 -0.400 14.410 0.400 ;
        RECT  14.410 -0.400 14.810 0.560 ;
        RECT  14.810 -0.400 16.900 0.400 ;
        RECT  16.900 -0.400 16.910 1.020 ;
        RECT  16.910 -0.400 17.310 1.220 ;
        RECT  17.310 -0.400 17.320 1.020 ;
        RECT  17.320 -0.400 18.160 0.400 ;
        RECT  18.160 -0.400 18.170 0.690 ;
        RECT  18.170 -0.400 18.570 0.890 ;
        RECT  18.570 -0.400 18.580 0.690 ;
        RECT  18.580 -0.400 19.680 0.400 ;
        RECT  19.680 -0.400 19.690 0.790 ;
        RECT  19.690 -0.400 20.090 0.990 ;
        RECT  20.090 -0.400 20.100 0.790 ;
        RECT  20.100 -0.400 21.210 0.400 ;
        RECT  21.210 -0.400 21.610 1.460 ;
        RECT  21.610 -0.400 21.780 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  21.260 2.030 21.500 3.730 ;
        RECT  21.250 2.030 21.260 2.430 ;
        RECT  18.650 3.490 21.260 3.730 ;
        RECT  18.410 1.390 18.650 3.730 ;
        RECT  18.070 1.390 18.410 1.630 ;
        RECT  17.710 2.890 18.410 3.290 ;
        RECT  16.820 2.050 18.170 2.450 ;
        RECT  17.670 1.230 18.070 1.630 ;
        RECT  16.670 1.500 16.820 3.210 ;
        RECT  16.580 1.500 16.670 3.370 ;
        RECT  16.090 1.500 16.580 1.740 ;
        RECT  16.270 2.970 16.580 3.370 ;
        RECT  15.400 2.100 16.300 2.500 ;
        RECT  15.230 2.970 16.270 3.210 ;
        RECT  15.690 1.050 16.090 1.740 ;
        RECT  14.060 1.050 15.690 1.290 ;
        RECT  13.500 2.180 15.400 2.420 ;
        RECT  15.070 2.970 15.230 3.370 ;
        RECT  14.830 2.970 15.070 3.730 ;
        RECT  13.770 3.490 14.830 3.730 ;
        RECT  13.530 3.490 13.770 4.070 ;
        RECT  12.000 0.860 13.680 1.100 ;
        RECT  13.460 1.380 13.500 2.420 ;
        RECT  13.260 1.380 13.460 3.090 ;
        RECT  13.040 1.380 13.260 1.780 ;
        RECT  13.220 2.180 13.260 3.090 ;
        RECT  13.040 2.850 13.220 3.090 ;
        RECT  11.480 1.380 13.040 1.620 ;
        RECT  12.800 2.850 13.040 3.310 ;
        RECT  12.740 2.170 12.980 2.570 ;
        RECT  11.330 3.070 12.800 3.310 ;
        RECT  11.820 2.170 12.740 2.410 ;
        RECT  11.760 0.670 12.000 1.100 ;
        RECT  11.580 1.860 11.820 2.410 ;
        RECT  10.790 0.670 11.760 0.910 ;
        RECT  11.380 1.860 11.580 2.100 ;
        RECT  11.080 1.190 11.480 1.620 ;
        RECT  10.930 3.070 11.330 3.470 ;
        RECT  10.800 2.280 11.100 2.680 ;
        RECT  10.660 2.270 10.800 2.680 ;
        RECT  10.660 0.670 10.790 1.630 ;
        RECT  10.550 0.670 10.660 3.270 ;
        RECT  10.420 1.390 10.550 3.270 ;
        RECT  9.320 1.390 10.420 1.650 ;
        RECT  9.140 3.030 10.420 3.270 ;
        RECT  8.860 2.230 10.140 2.640 ;
        RECT  9.160 1.240 9.320 1.650 ;
        RECT  9.000 3.550 9.240 4.130 ;
        RECT  9.000 0.670 9.160 1.650 ;
        RECT  8.920 0.670 9.000 1.640 ;
        RECT  6.580 3.550 9.000 3.790 ;
        RECT  8.860 0.670 8.920 1.070 ;
        RECT  8.620 1.930 8.860 3.270 ;
        RECT  8.500 1.930 8.620 2.170 ;
        RECT  7.100 3.030 8.620 3.270 ;
        RECT  8.260 0.930 8.500 2.170 ;
        RECT  7.930 2.450 8.340 2.690 ;
        RECT  7.690 1.400 7.930 2.690 ;
        RECT  5.960 1.400 7.690 1.640 ;
        RECT  6.860 2.180 7.100 3.270 ;
        RECT  6.840 2.180 6.860 2.580 ;
        RECT  6.560 2.850 6.580 4.350 ;
        RECT  6.340 1.990 6.560 4.350 ;
        RECT  6.320 1.990 6.340 3.090 ;
        RECT  4.440 4.110 6.340 4.350 ;
        RECT  6.090 1.990 6.320 2.390 ;
        RECT  5.820 3.360 6.060 3.760 ;
        RECT  5.810 0.990 5.960 1.640 ;
        RECT  5.810 3.360 5.820 3.600 ;
        RECT  5.570 0.990 5.810 3.600 ;
        RECT  5.560 0.990 5.570 1.390 ;
        RECT  4.860 3.130 5.260 3.620 ;
        RECT  4.680 0.860 5.080 1.290 ;
        RECT  2.390 3.130 4.860 3.370 ;
        RECT  2.380 0.860 4.680 1.100 ;
        RECT  4.200 3.670 4.440 4.350 ;
        RECT  3.130 3.670 4.200 3.910 ;
        RECT  2.380 1.380 4.040 1.620 ;
        RECT  2.890 3.670 3.130 4.110 ;
        RECT  2.380 2.540 3.090 2.780 ;
        RECT  0.570 3.870 2.890 4.110 ;
        RECT  1.980 0.670 2.380 1.100 ;
        RECT  2.140 1.380 2.380 2.780 ;
        RECT  2.110 2.540 2.140 2.780 ;
        RECT  1.870 2.540 2.110 3.590 ;
        RECT  1.650 3.350 1.870 3.590 ;
        RECT  0.490 1.240 0.570 1.640 ;
        RECT  0.490 2.930 0.570 4.110 ;
        RECT  0.330 1.240 0.490 4.110 ;
        RECT  0.250 1.240 0.330 3.330 ;
        RECT  0.170 1.240 0.250 1.640 ;
        RECT  0.170 2.930 0.250 3.330 ;
    END
END SDFFNSX4

MACRO SDFFNSX2
    CLASS CORE ;
    FOREIGN SDFFNSX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNSXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.800 1.830 7.060 2.090 ;
        RECT  7.060 1.840 7.460 2.400 ;
        RECT  7.460 1.840 7.470 2.320 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.280 2.010 3.760 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.470 1.460 1.870 2.270 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.150 2.750 15.190 3.150 ;
        RECT  15.030 0.670 15.190 0.910 ;
        RECT  15.190 0.670 15.370 3.150 ;
        RECT  15.370 0.670 15.430 3.160 ;
        RECT  15.430 2.390 15.640 3.160 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.040 1.270 16.150 1.530 ;
        RECT  16.150 1.260 16.590 1.540 ;
        RECT  16.590 0.700 16.710 1.680 ;
        RECT  16.590 3.130 16.750 4.110 ;
        RECT  16.710 0.700 16.750 1.840 ;
        RECT  16.750 0.700 16.990 4.110 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 1.760 4.700 2.160 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.700 2.100 1.170 2.660 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.210 5.440 ;
        RECT  0.210 4.480 0.610 5.440 ;
        RECT  0.610 4.640 3.370 5.440 ;
        RECT  3.370 4.110 3.610 5.440 ;
        RECT  3.610 4.640 6.700 5.440 ;
        RECT  6.700 4.480 7.100 5.440 ;
        RECT  7.100 4.640 8.220 5.440 ;
        RECT  8.220 4.310 8.230 5.440 ;
        RECT  8.230 4.190 8.630 5.440 ;
        RECT  8.630 4.310 8.640 5.440 ;
        RECT  8.640 4.640 9.620 5.440 ;
        RECT  9.620 3.880 9.630 5.440 ;
        RECT  9.630 3.680 10.030 5.440 ;
        RECT  10.030 3.880 10.040 5.440 ;
        RECT  10.040 4.640 12.120 5.440 ;
        RECT  12.120 4.010 12.360 5.440 ;
        RECT  12.360 4.640 13.670 5.440 ;
        RECT  13.670 4.480 14.070 5.440 ;
        RECT  14.070 4.640 15.820 5.440 ;
        RECT  15.820 4.290 15.830 5.440 ;
        RECT  15.830 4.090 16.230 5.440 ;
        RECT  16.230 4.290 16.240 5.440 ;
        RECT  16.240 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.190 0.400 ;
        RECT  1.190 -0.400 1.590 0.560 ;
        RECT  1.590 -0.400 3.260 0.400 ;
        RECT  3.260 -0.400 3.660 0.560 ;
        RECT  3.660 -0.400 6.890 0.400 ;
        RECT  6.890 -0.400 6.900 0.910 ;
        RECT  6.900 -0.400 7.300 1.030 ;
        RECT  7.300 -0.400 7.310 0.910 ;
        RECT  7.310 -0.400 9.320 0.400 ;
        RECT  9.320 -0.400 9.560 1.110 ;
        RECT  9.560 -0.400 12.100 0.400 ;
        RECT  12.100 -0.400 12.110 0.760 ;
        RECT  12.110 -0.400 12.510 0.960 ;
        RECT  12.510 -0.400 12.520 0.760 ;
        RECT  12.520 -0.400 13.880 0.400 ;
        RECT  13.880 -0.400 14.280 0.560 ;
        RECT  14.280 -0.400 15.820 0.400 ;
        RECT  15.820 -0.400 15.830 0.790 ;
        RECT  15.830 -0.400 16.230 0.990 ;
        RECT  16.230 -0.400 16.240 0.790 ;
        RECT  16.240 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.310 2.170 16.470 2.570 ;
        RECT  16.070 2.170 16.310 3.740 ;
        RECT  14.870 3.500 16.070 3.740 ;
        RECT  14.870 1.330 14.890 1.730 ;
        RECT  14.630 1.330 14.870 3.740 ;
        RECT  14.490 1.330 14.630 1.730 ;
        RECT  14.330 3.340 14.630 3.740 ;
        RECT  14.210 2.020 14.350 2.450 ;
        RECT  13.970 1.510 14.210 3.060 ;
        RECT  13.010 1.510 13.970 1.750 ;
        RECT  13.260 2.820 13.970 3.060 ;
        RECT  13.100 2.820 13.260 3.380 ;
        RECT  12.860 2.820 13.100 3.730 ;
        RECT  12.610 1.240 13.010 1.750 ;
        RECT  11.820 3.490 12.860 3.730 ;
        RECT  12.400 2.100 12.800 2.500 ;
        RECT  11.810 1.240 12.610 1.480 ;
        RECT  11.590 2.180 12.400 2.420 ;
        RECT  11.580 3.490 11.820 4.070 ;
        RECT  11.350 1.880 11.590 3.160 ;
        RECT  11.420 3.670 11.580 4.070 ;
        RECT  11.170 0.670 11.410 1.560 ;
        RECT  10.840 1.880 11.350 2.120 ;
        RECT  11.230 2.920 11.350 3.160 ;
        RECT  10.990 2.920 11.230 3.330 ;
        RECT  10.320 0.670 11.170 0.910 ;
        RECT  10.320 2.400 11.050 2.640 ;
        RECT  10.600 1.190 10.840 2.120 ;
        RECT  10.080 0.670 10.320 3.180 ;
        RECT  9.030 1.390 10.080 1.650 ;
        RECT  9.510 2.940 10.080 3.180 ;
        RECT  9.560 1.930 9.800 2.330 ;
        RECT  8.830 1.970 9.560 2.210 ;
        RECT  9.110 2.940 9.510 3.340 ;
        RECT  8.910 3.670 9.150 4.070 ;
        RECT  8.790 0.670 9.030 1.650 ;
        RECT  6.350 3.670 8.910 3.910 ;
        RECT  8.590 1.970 8.830 3.390 ;
        RECT  7.790 0.670 8.790 0.910 ;
        RECT  8.510 1.970 8.590 2.210 ;
        RECT  6.870 3.150 8.590 3.390 ;
        RECT  8.270 1.430 8.510 2.210 ;
        RECT  7.990 2.520 8.310 2.760 ;
        RECT  7.750 1.310 7.990 2.760 ;
        RECT  6.620 1.310 7.750 1.550 ;
        RECT  6.630 2.720 6.870 3.390 ;
        RECT  6.380 1.150 6.620 1.550 ;
        RECT  5.880 1.150 6.380 1.390 ;
        RECT  6.110 1.830 6.350 4.100 ;
        RECT  6.100 1.830 6.110 2.070 ;
        RECT  4.290 3.860 6.110 4.100 ;
        RECT  5.860 1.670 6.100 2.070 ;
        RECT  5.580 0.860 5.880 1.390 ;
        RECT  5.590 2.640 5.830 3.580 ;
        RECT  5.580 2.640 5.590 2.880 ;
        RECT  5.480 0.860 5.580 2.880 ;
        RECT  5.340 1.150 5.480 2.880 ;
        RECT  4.630 3.070 5.030 3.570 ;
        RECT  4.600 0.850 5.000 1.250 ;
        RECT  2.570 3.070 4.630 3.310 ;
        RECT  2.320 0.860 4.600 1.100 ;
        RECT  4.050 3.590 4.290 4.100 ;
        RECT  3.090 3.590 4.050 3.830 ;
        RECT  2.380 1.380 3.800 1.620 ;
        RECT  2.850 3.590 3.090 4.370 ;
        RECT  2.380 2.540 2.870 2.780 ;
        RECT  1.840 4.130 2.850 4.370 ;
        RECT  2.330 3.070 2.570 3.850 ;
        RECT  2.140 1.380 2.380 2.780 ;
        RECT  2.170 3.610 2.330 3.850 ;
        RECT  1.920 0.670 2.320 1.100 ;
        RECT  2.050 2.540 2.140 2.780 ;
        RECT  1.810 2.540 2.050 3.110 ;
        RECT  1.600 3.790 1.840 4.370 ;
        RECT  1.650 2.870 1.810 3.110 ;
        RECT  0.570 3.790 1.600 4.030 ;
        RECT  0.430 1.270 0.730 1.670 ;
        RECT  0.430 2.930 0.570 4.030 ;
        RECT  0.330 1.270 0.430 4.030 ;
        RECT  0.190 1.270 0.330 3.330 ;
        RECT  0.170 2.930 0.190 3.330 ;
    END
END SDFFNSX2

MACRO SDFFNSX1
    CLASS CORE ;
    FOREIGN SDFFNSX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNSXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  12.650 3.930 13.210 4.350 ;
        RECT  13.210 3.940 13.280 4.340 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.410 2.150 3.810 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.470 1.700 1.870 2.250 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.340 3.650 14.640 4.050 ;
        RECT  14.640 3.510 14.740 4.050 ;
        RECT  14.340 0.670 14.740 1.100 ;
        RECT  14.740 3.500 14.880 4.050 ;
        RECT  14.880 3.500 14.980 3.770 ;
        RECT  14.980 3.500 15.300 3.740 ;
        RECT  14.740 0.860 15.300 1.100 ;
        RECT  15.300 0.860 15.540 3.740 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.930 2.840 15.950 3.240 ;
        RECT  15.930 1.220 15.950 1.620 ;
        RECT  15.950 1.210 16.340 3.250 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.950 1.520 4.070 1.760 ;
        RECT  4.070 1.510 4.510 2.100 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.290 0.800 2.690 ;
        RECT  0.800 2.280 1.130 2.700 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.780 5.440 ;
        RECT  0.780 4.480 1.180 5.440 ;
        RECT  1.180 4.640 3.500 5.440 ;
        RECT  3.500 4.270 3.510 5.440 ;
        RECT  3.510 4.150 3.910 5.440 ;
        RECT  3.910 4.270 3.920 5.440 ;
        RECT  3.920 4.640 6.860 5.440 ;
        RECT  6.860 4.480 7.260 5.440 ;
        RECT  7.260 4.640 8.280 5.440 ;
        RECT  8.280 4.210 8.290 5.440 ;
        RECT  8.290 4.090 8.690 5.440 ;
        RECT  8.690 4.210 8.700 5.440 ;
        RECT  8.700 4.640 9.590 5.440 ;
        RECT  9.590 3.790 9.600 5.440 ;
        RECT  9.600 3.590 10.000 5.440 ;
        RECT  10.000 3.790 10.010 5.440 ;
        RECT  10.010 4.640 11.930 5.440 ;
        RECT  11.930 3.790 11.940 5.440 ;
        RECT  11.940 3.590 12.340 5.440 ;
        RECT  12.340 3.790 12.350 5.440 ;
        RECT  12.350 4.640 13.550 5.440 ;
        RECT  13.520 3.080 13.550 3.480 ;
        RECT  13.550 3.070 13.970 5.440 ;
        RECT  13.970 4.640 15.130 5.440 ;
        RECT  15.130 4.480 15.530 5.440 ;
        RECT  15.530 4.640 16.500 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.830 0.400 ;
        RECT  0.830 -0.400 1.230 0.560 ;
        RECT  1.230 -0.400 2.910 0.400 ;
        RECT  2.910 -0.400 3.310 0.560 ;
        RECT  3.310 -0.400 6.460 0.400 ;
        RECT  6.460 -0.400 6.470 0.880 ;
        RECT  6.470 -0.400 6.870 1.000 ;
        RECT  6.870 -0.400 6.880 0.880 ;
        RECT  6.880 -0.400 9.130 0.400 ;
        RECT  9.130 -0.400 9.370 0.950 ;
        RECT  9.370 -0.400 11.510 0.400 ;
        RECT  11.510 -0.400 11.910 0.560 ;
        RECT  11.910 -0.400 13.570 0.400 ;
        RECT  13.570 -0.400 13.580 0.670 ;
        RECT  13.580 -0.400 13.980 0.870 ;
        RECT  13.980 -0.400 13.990 0.670 ;
        RECT  13.990 -0.400 14.990 0.400 ;
        RECT  14.990 -0.400 15.540 0.620 ;
        RECT  15.540 -0.400 16.500 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.780 1.380 15.020 3.230 ;
        RECT  14.400 1.380 14.780 1.780 ;
        RECT  14.400 2.990 14.780 3.230 ;
        RECT  13.820 2.110 14.220 2.510 ;
        RECT  13.160 2.190 13.820 2.430 ;
        RECT  12.920 1.630 13.160 3.430 ;
        RECT  12.700 1.630 12.920 1.870 ;
        RECT  12.760 3.030 12.920 3.430 ;
        RECT  12.300 1.160 12.700 1.870 ;
        RECT  12.400 2.350 12.640 2.750 ;
        RECT  11.140 2.510 12.400 2.750 ;
        RECT  11.860 1.630 12.300 1.870 ;
        RECT  11.460 1.630 11.860 2.030 ;
        RECT  11.140 3.520 11.220 3.920 ;
        RECT  10.900 1.350 11.140 3.920 ;
        RECT  10.110 0.670 11.090 0.910 ;
        RECT  10.790 1.350 10.900 1.590 ;
        RECT  10.820 3.520 10.900 3.920 ;
        RECT  10.390 1.190 10.790 1.590 ;
        RECT  10.110 2.510 10.620 2.920 ;
        RECT  9.870 0.670 10.110 2.920 ;
        RECT  8.810 1.230 9.870 1.470 ;
        RECT  9.670 2.680 9.870 2.920 ;
        RECT  9.270 2.680 9.670 3.180 ;
        RECT  8.950 1.750 9.590 2.150 ;
        RECT  9.050 3.570 9.290 4.070 ;
        RECT  6.570 3.570 9.050 3.810 ;
        RECT  8.710 1.750 8.950 3.290 ;
        RECT  8.570 0.670 8.810 1.470 ;
        RECT  8.290 1.750 8.710 1.990 ;
        RECT  7.110 3.050 8.710 3.290 ;
        RECT  7.150 0.670 8.570 0.910 ;
        RECT  8.030 2.370 8.430 2.770 ;
        RECT  8.050 1.370 8.290 1.990 ;
        RECT  7.630 2.370 8.030 2.610 ;
        RECT  7.390 1.280 7.630 2.610 ;
        RECT  5.530 1.280 7.390 1.520 ;
        RECT  6.870 2.130 7.110 3.290 ;
        RECT  6.810 2.130 6.870 2.370 ;
        RECT  6.570 1.970 6.810 2.370 ;
        RECT  6.330 2.650 6.570 4.090 ;
        RECT  6.290 2.650 6.330 2.890 ;
        RECT  4.510 3.850 6.330 4.090 ;
        RECT  6.050 1.800 6.290 2.890 ;
        RECT  5.430 1.800 6.050 2.040 ;
        RECT  5.810 3.160 6.050 3.560 ;
        RECT  5.770 3.160 5.810 3.400 ;
        RECT  5.530 2.590 5.770 3.400 ;
        RECT  5.150 1.000 5.530 1.520 ;
        RECT  5.150 2.590 5.530 2.830 ;
        RECT  4.850 3.110 5.250 3.420 ;
        RECT  5.130 1.000 5.150 2.830 ;
        RECT  4.910 1.280 5.130 2.830 ;
        RECT  2.390 3.110 4.850 3.350 ;
        RECT  4.330 0.840 4.570 1.240 ;
        RECT  4.270 3.630 4.510 4.090 ;
        RECT  1.970 0.860 4.330 1.100 ;
        RECT  0.570 3.630 4.270 3.870 ;
        RECT  2.380 1.380 3.610 1.620 ;
        RECT  2.380 2.540 3.090 2.780 ;
        RECT  2.140 1.380 2.380 2.780 ;
        RECT  2.050 2.540 2.140 2.780 ;
        RECT  1.810 2.540 2.050 3.280 ;
        RECT  1.570 0.670 1.970 1.100 ;
        RECT  1.650 2.880 1.810 3.280 ;
        RECT  0.400 1.330 0.570 1.730 ;
        RECT  0.400 2.970 0.570 3.870 ;
        RECT  0.330 1.330 0.400 3.870 ;
        RECT  0.160 1.330 0.330 3.410 ;
    END
END SDFFNSX1

MACRO SDFFNRXL
    CLASS CORE ;
    FOREIGN SDFFNRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.820 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.160 2.320 3.170 2.690 ;
        RECT  3.170 2.060 3.570 2.690 ;
        RECT  3.570 2.320 3.580 2.690 ;
        RECT  3.580 2.390 3.760 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 1.820 1.870 2.280 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.800 2.390 6.930 2.650 ;
        RECT  6.930 2.390 7.060 3.190 ;
        RECT  7.060 2.400 7.170 3.190 ;
        RECT  7.170 2.940 7.370 3.190 ;
        RECT  7.370 2.950 7.610 3.190 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.960 0.720 15.970 1.100 ;
        RECT  15.830 3.690 16.230 4.090 ;
        RECT  15.970 0.710 16.370 1.100 ;
        RECT  16.230 3.690 16.760 3.930 ;
        RECT  16.370 0.860 16.760 1.100 ;
        RECT  16.760 0.860 17.000 3.930 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.330 1.390 17.360 1.820 ;
        RECT  17.330 3.040 17.370 3.460 ;
        RECT  17.360 1.390 17.370 2.090 ;
        RECT  17.370 1.390 17.610 3.460 ;
        RECT  17.610 1.830 17.620 2.090 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.940 1.640 3.950 2.100 ;
        RECT  3.950 1.610 4.410 2.100 ;
        RECT  4.410 1.640 4.420 2.100 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.740 2.310 1.170 2.730 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.360 5.440 ;
        RECT  0.360 4.480 0.760 5.440 ;
        RECT  0.760 4.640 3.390 5.440 ;
        RECT  3.390 4.310 3.400 5.440 ;
        RECT  3.400 4.190 3.800 5.440 ;
        RECT  3.800 4.310 3.810 5.440 ;
        RECT  3.810 4.640 6.940 5.440 ;
        RECT  6.940 4.480 7.340 5.440 ;
        RECT  7.340 4.640 10.410 5.440 ;
        RECT  10.410 4.110 11.390 5.440 ;
        RECT  11.390 4.640 13.740 5.440 ;
        RECT  13.740 4.180 13.750 5.440 ;
        RECT  13.750 3.980 14.150 5.440 ;
        RECT  14.150 4.180 14.160 5.440 ;
        RECT  14.160 4.640 16.640 5.440 ;
        RECT  16.640 4.480 17.040 5.440 ;
        RECT  17.040 4.640 17.820 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 2.910 0.400 ;
        RECT  2.910 -0.400 3.310 0.560 ;
        RECT  3.310 -0.400 6.610 0.400 ;
        RECT  6.610 -0.400 6.620 0.730 ;
        RECT  6.620 -0.400 7.020 0.850 ;
        RECT  7.020 -0.400 7.030 0.730 ;
        RECT  7.030 -0.400 8.710 0.400 ;
        RECT  8.710 -0.400 9.020 1.540 ;
        RECT  9.020 1.190 9.270 1.530 ;
        RECT  9.270 1.190 10.520 1.540 ;
        RECT  10.520 1.190 10.920 1.880 ;
        RECT  9.020 -0.400 13.200 0.400 ;
        RECT  13.200 -0.400 13.210 1.110 ;
        RECT  13.210 -0.400 13.610 1.310 ;
        RECT  13.610 -0.400 13.620 1.110 ;
        RECT  13.620 -0.400 15.080 0.400 ;
        RECT  15.080 -0.400 15.090 0.690 ;
        RECT  15.090 -0.400 15.490 0.890 ;
        RECT  15.490 -0.400 15.500 0.690 ;
        RECT  15.500 -0.400 17.050 0.400 ;
        RECT  17.050 -0.400 17.450 0.560 ;
        RECT  17.450 -0.400 17.820 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.240 1.450 16.480 3.150 ;
        RECT  15.970 1.450 16.240 1.690 ;
        RECT  16.090 2.910 16.240 3.150 ;
        RECT  15.850 2.910 16.090 3.340 ;
        RECT  15.540 1.970 15.840 2.370 ;
        RECT  15.430 1.590 15.540 3.590 ;
        RECT  15.300 1.590 15.430 3.750 ;
        RECT  14.610 1.590 15.300 1.830 ;
        RECT  15.030 3.350 15.300 3.750 ;
        RECT  14.620 2.110 15.020 2.510 ;
        RECT  13.190 2.270 14.620 2.510 ;
        RECT  14.210 1.130 14.610 1.830 ;
        RECT  13.310 1.590 14.210 1.830 ;
        RECT  12.910 1.590 13.310 1.940 ;
        RECT  12.950 2.270 13.190 3.780 ;
        RECT  12.120 2.270 12.950 2.510 ;
        RECT  12.930 3.540 12.950 3.780 ;
        RECT  12.530 3.540 12.930 3.940 ;
        RECT  12.270 2.790 12.670 3.100 ;
        RECT  11.580 0.670 12.560 0.910 ;
        RECT  11.580 2.790 12.270 3.030 ;
        RECT  11.880 1.330 12.120 2.510 ;
        RECT  11.340 0.670 11.580 3.030 ;
        RECT  9.290 0.670 11.340 0.910 ;
        RECT  11.100 2.760 11.340 3.030 ;
        RECT  10.860 2.760 11.100 3.450 ;
        RECT  9.530 2.230 11.060 2.470 ;
        RECT  10.290 2.870 10.530 3.830 ;
        RECT  10.140 3.590 10.290 3.830 ;
        RECT  9.900 3.590 10.140 4.370 ;
        RECT  7.850 4.130 9.900 4.370 ;
        RECT  9.290 1.820 9.530 3.690 ;
        RECT  8.440 1.820 9.290 2.060 ;
        RECT  9.190 3.450 9.290 3.690 ;
        RECT  8.790 3.450 9.190 3.850 ;
        RECT  8.370 2.340 9.010 2.580 ;
        RECT  8.200 1.110 8.440 2.060 ;
        RECT  8.130 2.340 8.370 3.850 ;
        RECT  8.070 1.110 8.200 1.890 ;
        RECT  7.920 2.340 8.130 2.580 ;
        RECT  6.570 1.650 8.070 1.890 ;
        RECT  7.520 2.170 7.920 2.580 ;
        RECT  7.610 3.940 7.850 4.370 ;
        RECT  7.540 0.770 7.770 1.010 ;
        RECT  6.530 3.940 7.610 4.180 ;
        RECT  7.300 0.770 7.540 1.370 ;
        RECT  5.530 1.130 7.300 1.370 ;
        RECT  6.170 1.650 6.570 2.110 ;
        RECT  6.440 2.930 6.530 4.350 ;
        RECT  6.290 2.390 6.440 4.350 ;
        RECT  6.200 2.390 6.290 3.170 ;
        RECT  4.320 4.110 6.290 4.350 ;
        RECT  5.890 2.390 6.200 2.630 ;
        RECT  5.850 3.520 6.010 3.760 ;
        RECT  5.650 1.710 5.890 2.630 ;
        RECT  5.610 2.910 5.850 3.760 ;
        RECT  5.530 1.710 5.650 2.110 ;
        RECT  5.370 2.910 5.610 3.150 ;
        RECT  5.250 0.950 5.530 1.370 ;
        RECT  5.250 2.630 5.370 3.150 ;
        RECT  5.130 0.950 5.250 3.150 ;
        RECT  4.930 3.430 5.170 3.840 ;
        RECT  5.010 0.950 5.130 2.870 ;
        RECT  4.850 3.430 4.930 3.670 ;
        RECT  4.610 3.150 4.850 3.670 ;
        RECT  4.250 0.860 4.650 1.330 ;
        RECT  2.410 3.150 4.610 3.390 ;
        RECT  4.080 3.670 4.320 4.350 ;
        RECT  2.160 0.860 4.250 1.100 ;
        RECT  0.570 3.670 4.080 3.910 ;
        RECT  2.380 1.420 3.610 1.660 ;
        RECT  2.380 2.580 2.850 2.820 ;
        RECT  2.140 1.420 2.380 2.820 ;
        RECT  1.920 0.670 2.160 1.100 ;
        RECT  1.990 2.580 2.140 2.820 ;
        RECT  1.750 2.580 1.990 3.270 ;
        RECT  1.570 0.670 1.920 0.910 ;
        RECT  0.400 1.360 0.570 1.760 ;
        RECT  0.400 3.010 0.570 3.910 ;
        RECT  0.330 1.360 0.400 3.910 ;
        RECT  0.170 1.360 0.330 3.410 ;
        RECT  0.160 1.360 0.170 3.330 ;
    END
END SDFFNRXL

MACRO SDFFNRX4
    CLASS CORE ;
    FOREIGN SDFFNRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNRXL ;
    SIZE 23.760 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.390 3.100 2.650 ;
        RECT  3.100 2.390 3.150 2.630 ;
        RECT  3.150 2.080 3.550 2.630 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 1.290 1.520 2.330 ;
        RECT  1.520 1.270 1.720 2.330 ;
        RECT  1.720 1.270 1.780 1.530 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.200 2.810 7.800 3.210 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  20.570 1.160 21.010 3.220 ;
        RECT  21.010 1.170 21.180 1.570 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.890 1.260 21.990 3.160 ;
        RECT  21.990 1.250 22.120 3.160 ;
        RECT  22.120 1.170 22.330 3.160 ;
        RECT  22.330 2.750 22.520 3.150 ;
        RECT  22.330 1.170 22.520 1.570 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.020 2.300 4.510 2.720 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.700 2.150 0.710 2.570 ;
        RECT  0.710 2.150 0.860 2.640 ;
        RECT  0.860 2.150 1.120 2.650 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.280 5.440 ;
        RECT  0.280 4.480 0.680 5.440 ;
        RECT  0.680 4.640 3.500 5.440 ;
        RECT  3.500 4.290 3.510 5.440 ;
        RECT  3.510 4.170 3.910 5.440 ;
        RECT  3.910 4.290 3.920 5.440 ;
        RECT  3.920 4.640 6.800 5.440 ;
        RECT  6.800 4.480 7.200 5.440 ;
        RECT  7.200 4.640 10.420 5.440 ;
        RECT  10.420 3.910 10.430 5.440 ;
        RECT  10.430 3.710 10.830 5.440 ;
        RECT  10.830 3.910 10.840 5.440 ;
        RECT  10.840 4.640 13.270 5.440 ;
        RECT  13.270 3.930 13.280 5.440 ;
        RECT  13.280 3.730 13.680 5.440 ;
        RECT  13.680 3.930 13.690 5.440 ;
        RECT  13.690 4.640 15.960 5.440 ;
        RECT  15.960 4.290 15.970 5.440 ;
        RECT  15.970 4.170 16.370 5.440 ;
        RECT  16.370 4.290 16.380 5.440 ;
        RECT  16.380 4.640 18.460 5.440 ;
        RECT  18.460 3.580 18.470 5.440 ;
        RECT  18.470 3.090 18.870 5.440 ;
        RECT  18.870 3.580 18.880 5.440 ;
        RECT  18.880 4.640 19.960 5.440 ;
        RECT  19.960 4.210 19.970 5.440 ;
        RECT  19.970 4.010 20.370 5.440 ;
        RECT  20.370 4.210 20.380 5.440 ;
        RECT  20.380 4.640 21.440 5.440 ;
        RECT  21.440 4.210 21.450 5.440 ;
        RECT  21.450 4.010 21.850 5.440 ;
        RECT  21.850 4.210 21.860 5.440 ;
        RECT  21.860 4.640 22.980 5.440 ;
        RECT  22.980 4.210 22.990 5.440 ;
        RECT  22.990 4.010 23.390 5.440 ;
        RECT  23.390 4.210 23.400 5.440 ;
        RECT  23.400 4.640 23.760 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.400 0.400 ;
        RECT  0.400 -0.400 0.800 0.560 ;
        RECT  0.800 -0.400 3.010 0.400 ;
        RECT  3.010 -0.400 3.410 0.560 ;
        RECT  3.410 -0.400 7.560 0.400 ;
        RECT  7.560 -0.400 8.540 1.290 ;
        RECT  8.540 -0.400 9.590 0.400 ;
        RECT  9.590 -0.400 9.600 0.890 ;
        RECT  9.600 -0.400 10.000 1.090 ;
        RECT  10.000 -0.400 10.010 0.890 ;
        RECT  10.010 -0.400 11.290 0.400 ;
        RECT  11.290 -0.400 11.300 1.110 ;
        RECT  11.300 -0.400 11.700 1.310 ;
        RECT  11.700 -0.400 11.710 1.110 ;
        RECT  11.710 -0.400 14.200 0.400 ;
        RECT  14.200 -0.400 14.600 0.560 ;
        RECT  14.600 -0.400 15.630 0.400 ;
        RECT  15.630 -0.400 15.640 0.710 ;
        RECT  15.640 -0.400 16.040 0.910 ;
        RECT  16.040 -0.400 16.050 0.710 ;
        RECT  16.050 -0.400 17.150 0.400 ;
        RECT  17.150 -0.400 17.160 0.700 ;
        RECT  17.160 -0.400 17.560 0.900 ;
        RECT  17.560 -0.400 17.570 0.700 ;
        RECT  17.570 -0.400 18.680 0.400 ;
        RECT  18.680 -0.400 18.690 0.710 ;
        RECT  18.690 -0.400 19.090 0.910 ;
        RECT  19.090 -0.400 19.100 0.710 ;
        RECT  19.100 -0.400 20.160 0.400 ;
        RECT  20.160 -0.400 20.170 0.690 ;
        RECT  20.170 -0.400 20.570 0.890 ;
        RECT  20.570 -0.400 20.580 0.690 ;
        RECT  20.580 -0.400 21.440 0.400 ;
        RECT  21.440 -0.400 21.450 0.690 ;
        RECT  21.450 -0.400 21.850 0.890 ;
        RECT  21.850 -0.400 21.860 0.690 ;
        RECT  21.860 -0.400 22.780 0.400 ;
        RECT  22.780 -0.400 22.790 0.690 ;
        RECT  22.790 -0.400 23.190 0.890 ;
        RECT  23.190 -0.400 23.200 0.690 ;
        RECT  23.200 -0.400 23.760 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  22.810 2.180 23.050 3.730 ;
        RECT  20.290 3.490 22.810 3.730 ;
        RECT  20.280 3.200 20.290 3.730 ;
        RECT  20.040 1.390 20.280 3.730 ;
        RECT  19.720 1.390 20.040 1.800 ;
        RECT  19.630 3.030 20.040 3.730 ;
        RECT  18.790 2.070 19.770 2.470 ;
        RECT  19.420 1.390 19.720 1.790 ;
        RECT  19.230 3.020 19.630 4.000 ;
        RECT  18.180 2.150 18.790 2.390 ;
        RECT  18.180 0.690 18.320 1.480 ;
        RECT  18.170 0.690 18.180 2.390 ;
        RECT  17.940 0.690 18.170 3.210 ;
        RECT  17.920 0.690 17.940 1.480 ;
        RECT  17.930 2.150 17.940 3.210 ;
        RECT  17.650 2.970 17.930 3.210 ;
        RECT  16.800 1.240 17.920 1.480 ;
        RECT  16.680 1.760 17.660 2.160 ;
        RECT  17.250 2.960 17.650 3.940 ;
        RECT  15.690 3.650 17.250 3.890 ;
        RECT  16.560 0.670 16.800 1.480 ;
        RECT  15.770 1.870 16.680 2.110 ;
        RECT  16.400 0.670 16.560 1.070 ;
        RECT  15.530 1.380 15.770 3.370 ;
        RECT  15.450 3.650 15.690 4.350 ;
        RECT  14.410 1.380 15.530 1.790 ;
        RECT  14.960 3.130 15.530 3.370 ;
        RECT  13.920 0.860 15.180 1.100 ;
        RECT  14.700 2.450 15.100 2.850 ;
        RECT  14.560 3.130 14.960 4.230 ;
        RECT  12.880 2.450 14.700 2.690 ;
        RECT  13.000 3.130 14.560 3.370 ;
        RECT  13.400 1.380 14.410 1.620 ;
        RECT  13.680 0.700 13.920 1.100 ;
        RECT  12.240 0.700 13.680 0.940 ;
        RECT  13.160 1.220 13.400 1.620 ;
        RECT  12.520 1.220 13.160 1.460 ;
        RECT  12.760 3.130 13.000 3.860 ;
        RECT  12.640 1.750 12.880 2.690 ;
        RECT  12.460 3.620 12.760 3.860 ;
        RECT  12.060 3.620 12.460 4.020 ;
        RECT  12.240 1.750 12.360 3.180 ;
        RECT  12.120 0.700 12.240 3.180 ;
        RECT  12.000 0.700 12.120 1.990 ;
        RECT  11.770 2.940 12.120 3.180 ;
        RECT  10.740 1.750 12.000 1.990 ;
        RECT  10.180 2.270 11.840 2.510 ;
        RECT  11.710 2.940 11.770 3.340 ;
        RECT  11.310 2.940 11.710 4.130 ;
        RECT  10.630 2.810 11.030 3.430 ;
        RECT  10.500 0.670 10.740 1.990 ;
        RECT  10.050 3.190 10.630 3.430 ;
        RECT  10.280 0.670 10.500 0.910 ;
        RECT  9.940 1.570 10.180 2.910 ;
        RECT  9.810 3.190 10.050 4.370 ;
        RECT  7.360 1.570 9.940 1.810 ;
        RECT  9.530 2.670 9.940 2.910 ;
        RECT  7.720 4.130 9.810 4.370 ;
        RECT  8.400 2.150 9.660 2.390 ;
        RECT  9.290 2.670 9.530 3.800 ;
        RECT  9.130 3.560 9.290 3.800 ;
        RECT  8.160 2.090 8.400 3.850 ;
        RECT  7.640 2.090 8.160 2.330 ;
        RECT  8.000 3.610 8.160 3.850 ;
        RECT  7.480 3.940 7.720 4.370 ;
        RECT  6.470 3.940 7.480 4.180 ;
        RECT  7.120 1.570 7.360 2.530 ;
        RECT  5.630 0.770 7.130 1.010 ;
        RECT  6.910 2.290 7.120 2.530 ;
        RECT  6.670 2.290 6.910 2.690 ;
        RECT  6.390 3.010 6.470 4.350 ;
        RECT  6.230 2.080 6.390 4.350 ;
        RECT  6.150 2.080 6.230 3.250 ;
        RECT  4.430 4.110 6.230 4.350 ;
        RECT  5.870 2.080 6.150 2.320 ;
        RECT  5.790 3.530 5.950 3.770 ;
        RECT  5.630 1.840 5.870 2.320 ;
        RECT  5.550 2.600 5.790 3.770 ;
        RECT  5.390 0.770 5.630 1.560 ;
        RECT  5.350 2.600 5.550 2.840 ;
        RECT  5.350 1.320 5.390 1.560 ;
        RECT  5.110 1.320 5.350 2.840 ;
        RECT  5.030 3.480 5.190 3.720 ;
        RECT  4.790 3.130 5.030 3.720 ;
        RECT  2.710 3.130 4.790 3.370 ;
        RECT  4.350 0.860 4.750 1.300 ;
        RECT  4.190 3.650 4.430 4.350 ;
        RECT  2.730 0.860 4.350 1.100 ;
        RECT  3.230 3.650 4.190 3.890 ;
        RECT  2.440 1.440 3.720 1.680 ;
        RECT  2.990 3.650 3.230 4.130 ;
        RECT  1.460 3.890 2.990 4.130 ;
        RECT  2.490 0.670 2.730 1.100 ;
        RECT  2.470 3.130 2.710 3.610 ;
        RECT  1.650 0.670 2.490 0.910 ;
        RECT  2.380 1.440 2.440 2.850 ;
        RECT  2.140 1.430 2.380 2.850 ;
        RECT  2.050 2.610 2.140 2.850 ;
        RECT  1.810 2.610 2.050 3.510 ;
        RECT  1.650 3.110 1.810 3.510 ;
        RECT  1.220 3.790 1.460 4.130 ;
        RECT  0.570 3.790 1.220 4.030 ;
        RECT  0.410 1.190 0.570 1.590 ;
        RECT  0.410 3.150 0.570 4.030 ;
        RECT  0.330 1.190 0.410 4.030 ;
        RECT  0.170 1.190 0.330 3.550 ;
    END
END SDFFNRX4

MACRO SDFFNRX2
    CLASS CORE ;
    FOREIGN SDFFNRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNRXL ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.770 2.020 2.840 2.640 ;
        RECT  2.840 2.020 3.100 2.650 ;
        RECT  3.100 2.020 3.170 2.420 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 1.280 1.520 2.300 ;
        RECT  1.520 1.270 1.720 2.300 ;
        RECT  1.720 1.270 1.780 1.530 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.800 2.950 6.810 3.210 ;
        RECT  6.810 2.710 7.060 3.210 ;
        RECT  7.060 2.710 7.560 3.110 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.040 2.920 17.120 3.320 ;
        RECT  17.120 2.610 17.130 3.320 ;
        RECT  17.040 0.730 17.130 1.710 ;
        RECT  17.130 0.730 17.370 3.320 ;
        RECT  17.370 2.390 17.440 3.320 ;
        RECT  17.370 0.730 17.440 1.710 ;
        RECT  17.440 2.390 17.620 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.570 0.730 18.590 1.710 ;
        RECT  18.590 0.730 18.680 1.820 ;
        RECT  18.570 3.170 18.690 4.150 ;
        RECT  18.680 0.730 18.690 2.090 ;
        RECT  18.690 0.730 18.930 4.150 ;
        RECT  18.930 0.730 18.940 2.090 ;
        RECT  18.930 3.170 18.970 4.150 ;
        RECT  18.940 0.730 18.970 1.960 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.940 1.510 4.420 2.100 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.060 0.770 2.460 ;
        RECT  0.770 1.820 1.130 2.470 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.340 5.440 ;
        RECT  0.340 4.480 0.740 5.440 ;
        RECT  0.740 4.640 3.660 5.440 ;
        RECT  3.660 4.290 3.670 5.440 ;
        RECT  3.670 4.090 4.070 5.440 ;
        RECT  4.070 4.290 4.080 5.440 ;
        RECT  4.080 4.640 6.650 5.440 ;
        RECT  6.650 4.480 7.050 5.440 ;
        RECT  7.050 4.640 9.950 5.440 ;
        RECT  9.950 4.010 11.490 5.440 ;
        RECT  11.490 4.640 13.510 5.440 ;
        RECT  13.510 4.110 13.520 5.440 ;
        RECT  13.520 3.910 13.920 5.440 ;
        RECT  13.920 4.110 13.930 5.440 ;
        RECT  13.930 4.640 15.470 5.440 ;
        RECT  15.470 3.500 15.480 5.440 ;
        RECT  15.480 3.300 15.880 5.440 ;
        RECT  15.880 3.500 15.890 5.440 ;
        RECT  15.890 4.640 17.800 5.440 ;
        RECT  17.800 4.320 17.810 5.440 ;
        RECT  17.810 4.120 18.210 5.440 ;
        RECT  18.210 4.320 18.220 5.440 ;
        RECT  18.220 4.640 19.140 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 2.920 0.400 ;
        RECT  2.920 -0.400 3.320 0.560 ;
        RECT  3.320 -0.400 7.510 0.400 ;
        RECT  7.510 -0.400 7.910 1.310 ;
        RECT  7.910 -0.400 9.000 0.400 ;
        RECT  9.000 -0.400 9.010 0.640 ;
        RECT  9.010 -0.400 9.410 0.930 ;
        RECT  9.410 -0.400 9.420 0.640 ;
        RECT  9.420 -0.400 10.700 0.400 ;
        RECT  10.700 -0.400 10.710 1.020 ;
        RECT  10.710 -0.400 11.110 1.140 ;
        RECT  11.110 -0.400 11.120 1.020 ;
        RECT  11.120 -0.400 13.790 0.400 ;
        RECT  13.790 -0.400 14.190 0.560 ;
        RECT  14.190 -0.400 15.360 0.400 ;
        RECT  15.360 -0.400 15.370 1.100 ;
        RECT  15.370 -0.400 15.770 1.300 ;
        RECT  15.770 -0.400 15.780 1.100 ;
        RECT  15.780 -0.400 17.800 0.400 ;
        RECT  17.800 -0.400 17.810 1.200 ;
        RECT  17.810 -0.400 18.210 1.690 ;
        RECT  18.210 -0.400 18.220 1.200 ;
        RECT  18.220 -0.400 19.140 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  18.290 2.200 18.320 2.600 ;
        RECT  18.050 2.200 18.290 3.840 ;
        RECT  16.760 3.600 18.050 3.840 ;
        RECT  16.520 1.080 16.760 3.840 ;
        RECT  16.190 1.080 16.520 1.480 ;
        RECT  16.300 2.920 16.520 3.320 ;
        RECT  15.290 1.950 16.240 2.350 ;
        RECT  15.050 1.580 15.290 3.020 ;
        RECT  15.010 1.580 15.050 1.820 ;
        RECT  14.660 2.780 15.050 3.020 ;
        RECT  14.610 0.940 15.010 1.820 ;
        RECT  14.370 2.100 14.770 2.500 ;
        RECT  14.260 2.780 14.660 3.900 ;
        RECT  13.740 1.580 14.610 1.820 ;
        RECT  13.060 2.260 14.370 2.500 ;
        RECT  13.420 2.780 14.260 3.020 ;
        RECT  13.340 1.580 13.740 1.980 ;
        RECT  12.820 2.090 13.060 3.490 ;
        RECT  12.310 2.090 12.820 2.330 ;
        RECT  12.780 3.250 12.820 3.490 ;
        RECT  12.380 3.250 12.780 3.650 ;
        RECT  11.760 0.670 12.720 0.910 ;
        RECT  11.840 2.610 12.540 2.850 ;
        RECT  12.070 1.230 12.310 2.330 ;
        RECT  11.760 2.610 11.840 3.270 ;
        RECT  11.520 0.670 11.760 3.270 ;
        RECT  10.230 1.420 11.520 1.710 ;
        RECT  10.940 3.030 11.520 3.270 ;
        RECT  11.000 1.990 11.240 2.390 ;
        RECT  9.490 1.990 11.000 2.230 ;
        RECT  10.540 3.030 10.940 3.430 ;
        RECT  10.020 2.510 10.600 2.750 ;
        RECT  10.100 1.310 10.230 1.710 ;
        RECT  10.090 0.880 10.100 1.710 ;
        RECT  9.830 0.670 10.090 1.710 ;
        RECT  9.780 2.510 10.020 3.730 ;
        RECT  9.690 0.670 9.830 0.910 ;
        RECT  9.580 3.490 9.780 3.730 ;
        RECT  9.340 3.490 9.580 4.310 ;
        RECT  9.250 1.590 9.490 3.190 ;
        RECT  7.570 4.070 9.340 4.310 ;
        RECT  8.830 1.590 9.250 1.830 ;
        RECT  9.020 2.950 9.250 3.190 ;
        RECT  8.780 2.950 9.020 3.790 ;
        RECT  8.730 2.110 8.970 2.510 ;
        RECT  8.430 1.270 8.830 1.830 ;
        RECT  8.620 3.390 8.780 3.790 ;
        RECT  8.090 2.110 8.730 2.350 ;
        RECT  6.570 1.590 8.430 1.830 ;
        RECT  7.850 2.110 8.090 3.790 ;
        RECT  7.550 2.110 7.850 2.350 ;
        RECT  7.330 3.940 7.570 4.310 ;
        RECT  6.350 3.940 7.330 4.180 ;
        RECT  6.830 0.670 7.230 1.090 ;
        RECT  5.530 0.670 6.830 0.910 ;
        RECT  6.330 1.590 6.570 2.270 ;
        RECT  6.110 2.560 6.350 4.250 ;
        RECT  6.170 1.870 6.330 2.270 ;
        RECT  5.890 2.560 6.110 2.800 ;
        RECT  4.650 4.010 6.110 4.250 ;
        RECT  5.650 1.480 5.890 2.800 ;
        RECT  5.590 3.090 5.830 3.490 ;
        RECT  5.530 1.480 5.650 1.880 ;
        RECT  5.370 3.090 5.590 3.330 ;
        RECT  5.240 0.670 5.530 1.200 ;
        RECT  5.240 2.160 5.370 3.330 ;
        RECT  5.210 0.670 5.240 3.330 ;
        RECT  5.130 0.800 5.210 3.330 ;
        RECT  5.000 0.800 5.130 2.400 ;
        RECT  4.610 2.760 4.850 3.170 ;
        RECT  4.250 0.860 4.650 1.220 ;
        RECT  4.410 3.450 4.650 4.250 ;
        RECT  2.770 2.930 4.610 3.170 ;
        RECT  3.290 3.450 4.410 3.690 ;
        RECT  2.570 0.860 4.250 1.100 ;
        RECT  2.380 1.380 3.610 1.620 ;
        RECT  3.050 3.450 3.290 4.220 ;
        RECT  1.280 3.980 3.050 4.220 ;
        RECT  2.530 2.930 2.770 3.330 ;
        RECT  2.330 0.670 2.570 1.100 ;
        RECT  2.250 1.380 2.380 2.050 ;
        RECT  1.570 0.670 2.330 0.910 ;
        RECT  2.140 1.380 2.250 3.700 ;
        RECT  2.010 1.810 2.140 3.700 ;
        RECT  1.850 2.810 2.010 3.700 ;
        RECT  1.710 2.810 1.850 3.210 ;
        RECT  1.040 3.080 1.280 4.220 ;
        RECT  0.570 3.080 1.040 3.320 ;
        RECT  0.400 2.920 0.570 3.320 ;
        RECT  0.400 1.310 0.490 1.710 ;
        RECT  0.160 1.310 0.400 3.320 ;
    END
END SDFFNRX2

MACRO SDFFNRX1
    CLASS CORE ;
    FOREIGN SDFFNRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNRXL ;
    SIZE 17.820 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.080 2.100 3.500 2.640 ;
        RECT  3.500 2.390 3.760 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.200 1.830 1.600 2.240 ;
        RECT  1.600 1.830 1.780 2.090 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.800 2.390 6.930 2.650 ;
        RECT  6.930 2.390 7.060 3.190 ;
        RECT  7.060 2.400 7.170 3.190 ;
        RECT  7.170 2.940 7.370 3.190 ;
        RECT  7.370 2.950 7.610 3.190 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.830 3.690 16.230 4.090 ;
        RECT  15.850 0.710 16.300 1.100 ;
        RECT  16.230 3.690 16.760 3.930 ;
        RECT  16.300 0.860 16.760 1.100 ;
        RECT  16.760 0.860 17.000 3.930 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.330 1.310 17.360 1.820 ;
        RECT  17.330 3.170 17.370 3.570 ;
        RECT  17.360 1.310 17.370 2.090 ;
        RECT  17.370 1.310 17.610 3.570 ;
        RECT  17.610 1.830 17.620 2.090 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.940 1.640 4.510 2.120 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.640 0.860 3.040 ;
        RECT  0.860 2.640 0.920 3.210 ;
        RECT  0.920 2.760 1.110 3.210 ;
        RECT  1.110 2.950 1.120 3.210 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.360 5.440 ;
        RECT  0.360 4.480 0.760 5.440 ;
        RECT  0.760 4.640 3.350 5.440 ;
        RECT  3.350 4.310 3.360 5.440 ;
        RECT  3.360 4.190 3.760 5.440 ;
        RECT  3.760 4.310 3.770 5.440 ;
        RECT  3.770 4.640 6.930 5.440 ;
        RECT  6.930 4.480 7.330 5.440 ;
        RECT  7.330 4.640 10.410 5.440 ;
        RECT  10.410 4.110 11.390 5.440 ;
        RECT  11.390 4.640 13.330 5.440 ;
        RECT  13.330 4.190 13.340 5.440 ;
        RECT  13.340 3.990 13.740 5.440 ;
        RECT  13.740 4.190 13.750 5.440 ;
        RECT  13.750 4.640 16.660 5.440 ;
        RECT  16.660 4.480 17.060 5.440 ;
        RECT  17.060 4.640 17.820 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.890 0.400 ;
        RECT  0.890 -0.400 1.290 0.560 ;
        RECT  1.290 -0.400 2.970 0.400 ;
        RECT  2.970 -0.400 3.370 0.560 ;
        RECT  3.370 -0.400 6.610 0.400 ;
        RECT  6.610 -0.400 6.620 0.730 ;
        RECT  6.620 -0.400 7.020 0.850 ;
        RECT  7.020 -0.400 7.030 0.730 ;
        RECT  7.030 -0.400 8.770 0.400 ;
        RECT  8.770 -0.400 9.010 1.530 ;
        RECT  9.010 1.190 9.270 1.530 ;
        RECT  9.270 1.190 10.520 1.540 ;
        RECT  10.520 1.190 10.920 1.880 ;
        RECT  9.010 -0.400 13.200 0.400 ;
        RECT  13.200 -0.400 13.210 1.110 ;
        RECT  13.210 -0.400 13.610 1.310 ;
        RECT  13.610 -0.400 13.620 1.110 ;
        RECT  13.620 -0.400 15.080 0.400 ;
        RECT  15.080 -0.400 15.090 0.690 ;
        RECT  15.090 -0.400 15.490 0.890 ;
        RECT  15.490 -0.400 15.500 0.690 ;
        RECT  15.500 -0.400 17.140 0.400 ;
        RECT  17.140 -0.400 17.540 0.560 ;
        RECT  17.540 -0.400 17.820 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.240 1.450 16.480 3.150 ;
        RECT  15.910 1.450 16.240 1.690 ;
        RECT  16.090 2.910 16.240 3.150 ;
        RECT  15.850 2.910 16.090 3.340 ;
        RECT  15.540 1.970 15.840 2.370 ;
        RECT  15.300 1.590 15.540 3.750 ;
        RECT  14.610 1.590 15.300 1.830 ;
        RECT  15.020 3.350 15.300 3.750 ;
        RECT  14.620 2.110 15.020 2.510 ;
        RECT  12.930 2.270 14.620 2.510 ;
        RECT  14.210 1.020 14.610 1.830 ;
        RECT  13.590 1.590 14.210 1.830 ;
        RECT  13.190 1.590 13.590 1.990 ;
        RECT  12.870 2.270 12.930 4.130 ;
        RECT  12.630 1.420 12.870 4.130 ;
        RECT  12.180 1.420 12.630 1.660 ;
        RECT  12.530 3.730 12.630 4.130 ;
        RECT  11.580 0.670 12.560 0.910 ;
        RECT  12.100 2.470 12.340 3.000 ;
        RECT  11.940 1.260 12.180 1.660 ;
        RECT  11.580 2.760 12.100 3.000 ;
        RECT  11.340 0.670 11.580 3.000 ;
        RECT  9.290 0.670 11.340 0.910 ;
        RECT  11.100 2.760 11.340 3.000 ;
        RECT  10.860 2.760 11.100 3.450 ;
        RECT  9.620 2.230 11.060 2.470 ;
        RECT  10.290 2.870 10.530 3.830 ;
        RECT  10.140 3.590 10.290 3.830 ;
        RECT  9.900 3.590 10.140 4.370 ;
        RECT  7.850 4.130 9.900 4.370 ;
        RECT  9.380 1.820 9.620 3.390 ;
        RECT  8.490 1.820 9.380 2.060 ;
        RECT  9.110 3.150 9.380 3.390 ;
        RECT  8.870 3.150 9.110 3.850 ;
        RECT  8.370 2.340 9.100 2.580 ;
        RECT  8.250 1.110 8.490 2.060 ;
        RECT  8.130 2.340 8.370 3.850 ;
        RECT  8.070 1.110 8.250 1.890 ;
        RECT  7.920 2.340 8.130 2.580 ;
        RECT  6.580 1.650 8.070 1.890 ;
        RECT  7.520 2.170 7.920 2.580 ;
        RECT  7.610 3.940 7.850 4.370 ;
        RECT  7.540 0.770 7.770 1.010 ;
        RECT  6.650 3.940 7.610 4.180 ;
        RECT  7.300 0.770 7.540 1.370 ;
        RECT  5.590 1.130 7.300 1.370 ;
        RECT  6.440 2.930 6.650 4.360 ;
        RECT  6.340 1.650 6.580 2.150 ;
        RECT  6.410 2.470 6.440 4.360 ;
        RECT  6.200 2.470 6.410 3.170 ;
        RECT  4.280 4.120 6.410 4.360 ;
        RECT  6.180 1.910 6.340 2.150 ;
        RECT  5.870 2.470 6.200 2.710 ;
        RECT  5.920 3.520 6.130 3.760 ;
        RECT  5.680 2.990 5.920 3.760 ;
        RECT  5.630 1.680 5.870 2.710 ;
        RECT  5.340 2.990 5.680 3.230 ;
        RECT  5.520 1.680 5.630 2.080 ;
        RECT  5.230 0.930 5.590 1.370 ;
        RECT  5.230 2.630 5.340 3.230 ;
        RECT  4.800 3.520 5.250 3.760 ;
        RECT  5.190 0.930 5.230 3.230 ;
        RECT  5.100 1.010 5.190 3.230 ;
        RECT  4.990 1.010 5.100 2.870 ;
        RECT  4.560 3.150 4.800 3.760 ;
        RECT  4.610 0.930 4.710 1.330 ;
        RECT  4.310 0.860 4.610 1.330 ;
        RECT  2.360 3.150 4.560 3.390 ;
        RECT  2.160 0.860 4.310 1.100 ;
        RECT  4.040 3.670 4.280 4.360 ;
        RECT  0.500 3.670 4.040 3.910 ;
        RECT  2.380 1.380 3.540 1.620 ;
        RECT  2.380 2.550 2.610 2.790 ;
        RECT  2.140 1.380 2.380 2.790 ;
        RECT  1.920 0.670 2.160 1.100 ;
        RECT  1.940 2.550 2.140 2.790 ;
        RECT  1.700 2.550 1.940 3.270 ;
        RECT  1.630 0.670 1.920 0.910 ;
        RECT  0.400 1.360 0.570 1.760 ;
        RECT  0.400 3.320 0.500 3.910 ;
        RECT  0.160 1.360 0.400 3.910 ;
    END
END SDFFNRX1

MACRO SDFFNXL
    CLASS CORE ;
    FOREIGN SDFFNXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.520 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.360 1.820 2.370 2.100 ;
        RECT  2.370 1.590 2.610 2.100 ;
        RECT  2.610 1.820 3.560 2.100 ;
        RECT  3.560 1.820 3.780 2.410 ;
        RECT  3.780 1.840 3.800 2.410 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.030 2.380 2.590 2.680 ;
        RECT  2.590 2.380 2.830 3.050 ;
        RECT  2.830 2.810 4.420 3.050 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.970 1.780 13.980 3.250 ;
        RECT  13.980 1.390 14.310 3.250 ;
        RECT  14.310 1.780 14.320 3.250 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.390 2.920 12.790 3.320 ;
        RECT  12.790 2.930 13.000 3.210 ;
        RECT  12.780 0.720 13.180 1.100 ;
        RECT  13.000 2.930 13.460 3.170 ;
        RECT  13.180 0.860 13.460 1.100 ;
        RECT  13.460 0.860 13.700 3.170 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.080 1.500 4.160 2.080 ;
        RECT  4.160 1.500 4.420 2.090 ;
        RECT  4.420 1.500 4.530 2.080 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.730 2.170 0.860 2.640 ;
        RECT  0.860 2.170 1.120 2.650 ;
        RECT  1.120 2.170 1.200 2.640 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.750 5.440 ;
        RECT  0.750 4.480 1.150 5.440 ;
        RECT  1.150 4.640 3.710 5.440 ;
        RECT  3.710 4.480 4.110 5.440 ;
        RECT  4.110 4.640 9.130 5.440 ;
        RECT  9.130 4.480 9.530 5.440 ;
        RECT  9.530 4.640 11.580 5.440 ;
        RECT  11.580 4.480 11.980 5.440 ;
        RECT  11.980 4.640 13.180 5.440 ;
        RECT  13.180 4.480 13.580 5.440 ;
        RECT  13.580 4.640 14.520 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 2.970 0.400 ;
        RECT  2.970 -0.400 3.370 0.560 ;
        RECT  3.370 -0.400 6.700 0.400 ;
        RECT  6.700 -0.400 6.710 1.060 ;
        RECT  6.710 -0.400 7.110 1.180 ;
        RECT  7.110 -0.400 7.120 1.060 ;
        RECT  7.120 -0.400 9.290 0.400 ;
        RECT  9.290 -0.400 9.300 1.380 ;
        RECT  9.300 -0.400 9.700 1.500 ;
        RECT  9.700 -0.400 9.710 1.380 ;
        RECT  9.710 -0.400 11.890 0.400 ;
        RECT  11.890 -0.400 11.900 0.880 ;
        RECT  11.900 -0.400 12.300 1.080 ;
        RECT  12.300 -0.400 12.310 0.880 ;
        RECT  12.310 -0.400 13.730 0.400 ;
        RECT  13.730 -0.400 14.130 0.560 ;
        RECT  14.130 -0.400 14.520 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.940 1.460 13.180 2.640 ;
        RECT  12.780 1.460 12.940 1.700 ;
        RECT  11.740 2.400 12.940 2.640 ;
        RECT  12.450 3.800 12.850 4.200 ;
        RECT  12.100 1.660 12.500 2.110 ;
        RECT  11.700 3.800 12.450 4.040 ;
        RECT  11.020 1.660 12.100 1.900 ;
        RECT  11.700 2.310 11.740 2.710 ;
        RECT  11.460 2.310 11.700 4.040 ;
        RECT  11.340 2.310 11.460 2.710 ;
        RECT  10.240 0.760 11.250 1.000 ;
        RECT  10.780 1.280 11.020 4.220 ;
        RECT  10.520 1.280 10.780 1.680 ;
        RECT  10.470 3.820 10.780 4.220 ;
        RECT  10.240 2.610 10.470 3.010 ;
        RECT  10.190 0.760 10.240 3.010 ;
        RECT  10.000 0.760 10.190 4.180 ;
        RECT  8.820 1.800 10.000 2.040 ;
        RECT  9.950 2.770 10.000 4.180 ;
        RECT  8.850 3.940 9.950 4.180 ;
        RECT  9.430 2.320 9.670 3.660 ;
        RECT  8.330 3.420 9.430 3.660 ;
        RECT  8.610 3.940 8.850 4.370 ;
        RECT  8.650 1.170 8.820 2.040 ;
        RECT  8.650 2.740 8.730 3.140 ;
        RECT  8.420 1.170 8.650 3.140 ;
        RECT  6.760 4.130 8.610 4.370 ;
        RECT  8.410 1.250 8.420 3.140 ;
        RECT  8.330 2.740 8.410 3.140 ;
        RECT  8.090 3.420 8.330 3.850 ;
        RECT  7.500 3.610 8.090 3.850 ;
        RECT  7.670 1.010 7.910 2.390 ;
        RECT  7.500 2.150 7.670 2.390 ;
        RECT  7.240 2.150 7.500 3.850 ;
        RECT  6.480 1.510 7.390 1.750 ;
        RECT  6.860 2.150 7.240 2.550 ;
        RECT  6.580 2.890 6.760 4.370 ;
        RECT  6.520 2.350 6.580 4.370 ;
        RECT  6.340 2.350 6.520 3.130 ;
        RECT  6.120 3.930 6.520 4.370 ;
        RECT  6.240 1.500 6.480 1.750 ;
        RECT  5.570 2.350 6.340 2.590 ;
        RECT  5.770 1.500 6.240 1.740 ;
        RECT  5.900 3.410 6.200 3.650 ;
        RECT  5.660 2.870 5.900 3.650 ;
        RECT  5.370 0.860 5.770 1.740 ;
        RECT  5.310 3.930 5.710 4.330 ;
        RECT  5.050 2.870 5.660 3.110 ;
        RECT  5.330 2.020 5.570 2.590 ;
        RECT  2.470 3.390 5.380 3.630 ;
        RECT  5.050 1.500 5.370 1.740 ;
        RECT  4.940 3.930 5.310 4.170 ;
        RECT  4.810 1.500 5.050 3.110 ;
        RECT  4.700 3.910 4.940 4.170 ;
        RECT  4.490 0.820 4.890 1.220 ;
        RECT  2.710 3.910 4.700 4.150 ;
        RECT  1.980 0.860 4.490 1.100 ;
        RECT  2.470 3.910 2.710 4.360 ;
        RECT  1.670 4.120 2.470 4.360 ;
        RECT  1.950 2.960 2.190 3.840 ;
        RECT  1.800 1.470 2.040 1.870 ;
        RECT  1.580 0.670 1.980 1.100 ;
        RECT  1.760 2.960 1.950 3.200 ;
        RECT  1.760 1.630 1.800 1.870 ;
        RECT  1.520 1.630 1.760 3.200 ;
        RECT  1.430 3.540 1.670 4.360 ;
        RECT  0.570 3.540 1.430 3.780 ;
        RECT  0.410 1.310 0.570 1.710 ;
        RECT  0.410 2.930 0.570 3.780 ;
        RECT  0.330 1.310 0.410 3.780 ;
        RECT  0.170 1.310 0.330 3.330 ;
    END
END SDFFNXL

MACRO SDFFNX4
    CLASS CORE ;
    FOREIGN SDFFNX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNXL ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.950 2.870 3.210 ;
        RECT  2.870 2.710 2.880 3.210 ;
        RECT  2.880 2.540 3.100 3.210 ;
        RECT  3.100 2.540 3.280 3.200 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.990 2.220 2.360 2.660 ;
        RECT  2.360 2.020 2.610 2.660 ;
        RECT  2.610 2.020 3.560 2.260 ;
        RECT  3.560 2.020 3.800 2.820 ;
        RECT  3.800 2.580 3.950 2.820 ;
        RECT  3.950 2.580 4.350 2.980 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.930 1.820 17.940 3.220 ;
        RECT  17.940 1.820 17.950 3.270 ;
        RECT  17.950 1.390 18.340 3.270 ;
        RECT  18.340 1.390 18.350 3.220 ;
        RECT  18.350 1.820 18.370 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.440 2.870 16.610 3.270 ;
        RECT  16.610 1.390 17.010 3.270 ;
        RECT  17.010 1.820 17.050 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.070 1.510 4.510 2.100 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.710 1.920 0.860 2.640 ;
        RECT  0.860 1.920 1.120 2.650 ;
        RECT  1.120 1.920 1.180 2.640 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 4.480 1.390 5.440 ;
        RECT  1.390 4.640 6.930 5.440 ;
        RECT  6.930 4.480 7.330 5.440 ;
        RECT  7.330 4.640 9.430 5.440 ;
        RECT  9.430 4.480 9.830 5.440 ;
        RECT  9.830 4.640 11.860 5.440 ;
        RECT  11.860 4.140 12.260 5.440 ;
        RECT  12.260 4.640 14.200 5.440 ;
        RECT  14.200 4.140 14.600 5.440 ;
        RECT  14.600 4.640 15.710 5.440 ;
        RECT  15.710 4.270 15.720 5.440 ;
        RECT  15.720 4.070 16.120 5.440 ;
        RECT  16.120 4.270 16.130 5.440 ;
        RECT  16.130 4.640 17.170 5.440 ;
        RECT  17.170 4.270 17.180 5.440 ;
        RECT  17.180 4.070 17.580 5.440 ;
        RECT  17.580 4.270 17.590 5.440 ;
        RECT  17.590 4.640 18.560 5.440 ;
        RECT  18.560 4.270 18.570 5.440 ;
        RECT  18.570 4.070 18.970 5.440 ;
        RECT  18.970 4.270 18.980 5.440 ;
        RECT  18.980 4.640 19.140 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.930 0.400 ;
        RECT  0.930 -0.400 1.330 1.040 ;
        RECT  1.330 -0.400 3.010 0.400 ;
        RECT  3.010 -0.400 3.410 0.560 ;
        RECT  3.410 -0.400 6.680 0.400 ;
        RECT  6.680 -0.400 7.080 1.310 ;
        RECT  7.080 -0.400 9.530 0.400 ;
        RECT  9.530 -0.400 9.930 1.400 ;
        RECT  9.930 -0.400 11.950 0.400 ;
        RECT  11.950 -0.400 12.350 1.310 ;
        RECT  12.350 -0.400 14.480 0.400 ;
        RECT  14.480 -0.400 14.880 0.560 ;
        RECT  14.880 -0.400 15.990 0.400 ;
        RECT  15.990 -0.400 16.390 1.110 ;
        RECT  16.390 -0.400 17.270 0.400 ;
        RECT  17.270 -0.400 17.280 0.910 ;
        RECT  17.280 -0.400 17.680 1.110 ;
        RECT  17.680 -0.400 17.690 0.910 ;
        RECT  17.690 -0.400 18.560 0.400 ;
        RECT  18.560 -0.400 18.570 0.910 ;
        RECT  18.570 -0.400 18.970 1.110 ;
        RECT  18.970 -0.400 18.980 0.910 ;
        RECT  18.980 -0.400 19.140 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  18.610 2.190 18.850 3.790 ;
        RECT  16.200 3.550 18.610 3.790 ;
        RECT  15.960 1.390 16.200 3.790 ;
        RECT  15.670 1.390 15.960 1.630 ;
        RECT  14.920 3.390 15.960 3.790 ;
        RECT  15.480 2.260 15.720 3.050 ;
        RECT  15.270 1.100 15.670 1.630 ;
        RECT  14.410 2.810 15.480 3.050 ;
        RECT  14.890 1.390 15.270 1.630 ;
        RECT  14.650 1.390 14.890 2.520 ;
        RECT  14.170 0.990 14.410 3.860 ;
        RECT  12.890 0.990 14.170 1.230 ;
        RECT  13.480 3.620 14.170 3.860 ;
        RECT  13.560 1.510 13.800 2.910 ;
        RECT  13.250 2.670 13.560 2.910 ;
        RECT  13.080 3.620 13.480 4.020 ;
        RECT  13.090 2.670 13.250 3.070 ;
        RECT  12.850 2.670 13.090 3.340 ;
        RECT  11.080 3.620 13.080 3.860 ;
        RECT  12.650 0.990 12.890 1.830 ;
        RECT  10.960 3.100 12.850 3.340 ;
        RECT  11.150 1.590 12.650 1.830 ;
        RECT  11.730 2.110 12.130 2.510 ;
        RECT  10.180 2.110 11.730 2.350 ;
        RECT  10.750 1.240 11.150 1.830 ;
        RECT  10.680 3.620 11.080 4.020 ;
        RECT  10.560 2.640 10.960 3.340 ;
        RECT  10.710 1.320 10.750 1.830 ;
        RECT  9.030 3.100 10.560 3.340 ;
        RECT  10.100 1.920 10.180 2.630 ;
        RECT  9.770 1.680 10.100 2.630 ;
        RECT  9.250 1.680 9.770 1.920 ;
        RECT  9.010 0.760 9.250 1.920 ;
        RECT  8.730 3.030 9.030 3.430 ;
        RECT  7.840 0.760 9.010 1.000 ;
        RECT  8.490 1.280 8.730 4.180 ;
        RECT  8.330 1.280 8.490 1.680 ;
        RECT  6.550 3.940 8.490 4.180 ;
        RECT  7.840 3.420 8.150 3.660 ;
        RECT  7.600 0.760 7.840 3.660 ;
        RECT  7.440 1.100 7.600 1.500 ;
        RECT  7.190 2.660 7.600 2.900 ;
        RECT  6.920 1.830 7.320 2.180 ;
        RECT  6.790 2.580 7.190 2.980 ;
        RECT  6.070 1.830 6.920 2.070 ;
        RECT  6.510 3.940 6.550 4.240 ;
        RECT  6.270 2.350 6.510 4.240 ;
        RECT  5.540 2.350 6.270 2.590 ;
        RECT  6.000 4.000 6.270 4.240 ;
        RECT  5.830 1.420 6.070 2.070 ;
        RECT  5.750 2.880 5.990 3.680 ;
        RECT  5.710 1.420 5.830 1.660 ;
        RECT  5.020 2.880 5.750 3.120 ;
        RECT  5.310 0.690 5.710 1.660 ;
        RECT  5.150 4.060 5.550 4.370 ;
        RECT  5.300 1.940 5.540 2.590 ;
        RECT  5.020 1.420 5.310 1.660 ;
        RECT  3.800 3.400 5.310 3.640 ;
        RECT  1.910 4.060 5.150 4.300 ;
        RECT  4.780 1.420 5.020 3.120 ;
        RECT  4.430 0.720 4.830 1.120 ;
        RECT  3.930 0.880 4.430 1.120 ;
        RECT  3.690 0.880 3.930 1.220 ;
        RECT  2.070 1.500 3.800 1.740 ;
        RECT  3.560 3.400 3.800 3.780 ;
        RECT  2.070 0.980 3.690 1.220 ;
        RECT  2.470 3.540 3.560 3.780 ;
        RECT  1.910 2.940 2.480 3.180 ;
        RECT  1.670 0.750 2.070 1.220 ;
        RECT  1.720 1.500 2.070 1.910 ;
        RECT  1.720 2.940 1.910 3.260 ;
        RECT  1.670 3.840 1.910 4.300 ;
        RECT  1.480 1.500 1.720 3.260 ;
        RECT  0.570 3.840 1.670 4.080 ;
        RECT  0.430 1.200 0.570 1.600 ;
        RECT  0.430 3.110 0.570 4.090 ;
        RECT  0.190 1.200 0.430 4.090 ;
        RECT  0.170 1.200 0.190 1.600 ;
        RECT  0.170 3.110 0.190 4.090 ;
    END
END SDFFNX4

MACRO SDFFNX2
    CLASS CORE ;
    FOREIGN SDFFNX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.360 1.820 2.370 2.100 ;
        RECT  2.370 1.590 2.610 2.100 ;
        RECT  2.610 1.820 3.530 2.100 ;
        RECT  3.530 1.820 3.770 2.410 ;
        RECT  3.770 1.820 3.780 2.100 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.000 2.390 2.590 2.660 ;
        RECT  2.590 2.390 2.830 3.050 ;
        RECT  2.830 2.810 4.290 3.050 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.530 3.130 16.610 4.110 ;
        RECT  16.450 0.730 16.610 1.710 ;
        RECT  16.610 0.730 16.770 4.110 ;
        RECT  16.770 0.730 16.850 4.100 ;
        RECT  16.850 2.390 16.960 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.650 3.130 15.050 3.530 ;
        RECT  14.700 0.690 15.110 1.100 ;
        RECT  15.050 3.130 15.480 3.370 ;
        RECT  15.110 0.860 15.480 1.100 ;
        RECT  15.480 0.860 15.720 3.370 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 1.560 4.510 2.090 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.730 2.170 0.860 2.640 ;
        RECT  0.860 2.170 1.120 2.650 ;
        RECT  1.120 2.170 1.180 2.640 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.730 5.440 ;
        RECT  0.730 4.480 1.130 5.440 ;
        RECT  1.130 4.640 3.640 5.440 ;
        RECT  3.640 4.480 4.040 5.440 ;
        RECT  4.040 4.640 8.950 5.440 ;
        RECT  8.950 4.480 9.350 5.440 ;
        RECT  9.350 4.640 11.500 5.440 ;
        RECT  11.500 4.480 11.900 5.440 ;
        RECT  11.900 4.640 13.740 5.440 ;
        RECT  13.740 4.480 14.140 5.440 ;
        RECT  14.140 4.640 15.520 5.440 ;
        RECT  15.520 4.480 15.920 5.440 ;
        RECT  15.920 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.300 0.400 ;
        RECT  0.300 -0.400 0.700 0.560 ;
        RECT  0.700 -0.400 2.890 0.400 ;
        RECT  2.890 -0.400 3.290 0.560 ;
        RECT  3.290 -0.400 6.670 0.400 ;
        RECT  6.670 -0.400 6.680 1.020 ;
        RECT  6.680 -0.400 7.080 1.220 ;
        RECT  7.080 -0.400 7.090 1.020 ;
        RECT  7.090 -0.400 9.290 0.400 ;
        RECT  9.290 -0.400 9.300 1.200 ;
        RECT  9.300 -0.400 9.700 1.400 ;
        RECT  9.700 -0.400 9.710 1.200 ;
        RECT  9.710 -0.400 11.740 0.400 ;
        RECT  11.740 -0.400 12.140 1.400 ;
        RECT  12.140 -0.400 13.920 0.400 ;
        RECT  13.920 -0.400 13.930 0.790 ;
        RECT  13.930 -0.400 14.330 0.990 ;
        RECT  14.330 -0.400 14.340 0.790 ;
        RECT  14.340 -0.400 15.630 0.400 ;
        RECT  15.630 -0.400 16.030 0.560 ;
        RECT  16.030 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.000 2.170 16.240 4.090 ;
        RECT  15.050 3.850 16.000 4.090 ;
        RECT  14.970 1.380 15.070 1.780 ;
        RECT  14.650 3.850 15.050 4.320 ;
        RECT  14.730 1.380 14.970 2.850 ;
        RECT  14.370 2.610 14.730 2.850 ;
        RECT  14.370 3.850 14.650 4.090 ;
        RECT  14.250 1.600 14.490 2.320 ;
        RECT  14.130 2.610 14.370 4.090 ;
        RECT  13.250 1.600 14.250 1.840 ;
        RECT  13.770 2.610 14.130 2.850 ;
        RECT  13.530 2.180 13.770 2.850 ;
        RECT  13.010 1.600 13.250 3.650 ;
        RECT  12.990 1.600 13.010 1.920 ;
        RECT  12.640 3.410 13.010 3.650 ;
        RECT  12.590 1.100 12.990 1.920 ;
        RECT  12.490 2.410 12.730 2.860 ;
        RECT  12.240 3.410 12.640 3.810 ;
        RECT  10.920 1.680 12.590 1.920 ;
        RECT  10.380 2.620 12.490 2.860 ;
        RECT  10.620 3.520 12.240 3.760 ;
        RECT  10.680 1.240 10.920 1.920 ;
        RECT  10.520 1.240 10.680 1.640 ;
        RECT  10.220 3.520 10.620 3.920 ;
        RECT  10.220 2.620 10.380 3.240 ;
        RECT  9.980 1.790 10.220 3.240 ;
        RECT  8.740 1.790 9.980 2.030 ;
        RECT  9.610 3.000 9.980 3.240 ;
        RECT  9.240 2.320 9.640 2.720 ;
        RECT  9.370 3.000 9.610 4.180 ;
        RECT  8.660 3.940 9.370 4.180 ;
        RECT  9.080 2.480 9.240 2.720 ;
        RECT  8.840 2.480 9.080 3.660 ;
        RECT  8.140 3.420 8.840 3.660 ;
        RECT  8.740 1.080 8.820 1.320 ;
        RECT  8.500 1.080 8.740 2.030 ;
        RECT  8.420 3.940 8.660 4.370 ;
        RECT  8.500 2.740 8.560 3.140 ;
        RECT  8.260 1.080 8.500 3.140 ;
        RECT  6.730 4.130 8.420 4.370 ;
        RECT  8.160 2.740 8.260 3.140 ;
        RECT  7.740 3.420 8.140 3.800 ;
        RECT  7.740 0.910 7.900 1.310 ;
        RECT  7.500 0.910 7.740 3.800 ;
        RECT  6.640 2.290 7.500 2.530 ;
        RECT  6.820 1.500 7.220 1.810 ;
        RECT  5.710 1.500 6.820 1.740 ;
        RECT  6.490 2.880 6.730 4.370 ;
        RECT  6.360 2.880 6.490 3.120 ;
        RECT  6.180 3.920 6.490 4.370 ;
        RECT  6.120 2.350 6.360 3.120 ;
        RECT  5.840 3.390 6.200 3.630 ;
        RECT  6.100 3.930 6.180 4.370 ;
        RECT  5.540 2.350 6.120 2.590 ;
        RECT  5.600 2.870 5.840 3.630 ;
        RECT  5.680 3.930 5.760 4.330 ;
        RECT  5.310 1.050 5.710 1.740 ;
        RECT  5.360 3.920 5.680 4.330 ;
        RECT  5.020 2.870 5.600 3.110 ;
        RECT  5.300 2.020 5.540 2.590 ;
        RECT  2.900 3.920 5.360 4.160 ;
        RECT  5.240 3.390 5.320 3.630 ;
        RECT  5.020 1.500 5.310 1.740 ;
        RECT  4.920 3.390 5.240 3.640 ;
        RECT  4.780 1.500 5.020 3.110 ;
        RECT  2.410 3.400 4.920 3.640 ;
        RECT  4.430 0.830 4.830 1.230 ;
        RECT  1.950 0.860 4.430 1.100 ;
        RECT  2.660 3.920 2.900 4.360 ;
        RECT  1.630 4.120 2.660 4.360 ;
        RECT  1.890 2.960 2.130 3.840 ;
        RECT  1.770 1.470 2.010 1.870 ;
        RECT  1.550 0.670 1.950 1.100 ;
        RECT  1.720 2.960 1.890 3.200 ;
        RECT  1.720 1.630 1.770 1.870 ;
        RECT  1.480 1.630 1.720 3.200 ;
        RECT  1.390 3.860 1.630 4.360 ;
        RECT  0.570 3.860 1.390 4.100 ;
        RECT  0.450 1.310 0.570 1.710 ;
        RECT  0.450 3.000 0.570 4.100 ;
        RECT  0.330 1.310 0.450 4.100 ;
        RECT  0.210 1.310 0.330 3.400 ;
        RECT  0.170 1.310 0.210 1.710 ;
        RECT  0.170 3.000 0.210 3.400 ;
    END
END SDFFNX2

MACRO SDFFNX1
    CLASS CORE ;
    FOREIGN SDFFNX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFNXL ;
    SIZE 14.520 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.390 1.820 2.400 2.100 ;
        RECT  2.400 1.590 2.640 2.100 ;
        RECT  2.640 1.820 3.560 2.100 ;
        RECT  3.560 1.820 3.800 2.410 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.000 2.390 2.590 2.660 ;
        RECT  2.590 2.390 2.830 2.930 ;
        RECT  2.830 2.690 3.920 2.930 ;
        RECT  3.920 2.690 4.340 3.050 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.950 1.320 13.970 1.720 ;
        RECT  13.970 1.320 14.350 3.410 ;
        RECT  14.350 1.430 14.360 3.410 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.400 3.130 12.800 3.530 ;
        RECT  12.510 0.690 13.080 1.100 ;
        RECT  12.800 3.130 13.430 3.370 ;
        RECT  13.080 0.860 13.430 1.100 ;
        RECT  13.430 0.860 13.670 3.370 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.130 1.570 4.520 2.210 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.730 2.170 1.110 2.650 ;
        RECT  1.110 2.390 1.120 2.650 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.730 5.440 ;
        RECT  0.730 4.480 1.130 5.440 ;
        RECT  1.130 4.640 3.740 5.440 ;
        RECT  3.740 4.480 4.140 5.440 ;
        RECT  4.140 4.640 9.130 5.440 ;
        RECT  9.130 4.480 9.530 5.440 ;
        RECT  9.530 4.640 11.590 5.440 ;
        RECT  11.590 4.480 11.990 5.440 ;
        RECT  11.990 4.640 13.190 5.440 ;
        RECT  13.190 4.480 13.590 5.440 ;
        RECT  13.590 4.640 14.520 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 2.950 0.400 ;
        RECT  2.950 -0.400 3.350 0.560 ;
        RECT  3.350 -0.400 6.730 0.400 ;
        RECT  6.730 -0.400 6.740 1.030 ;
        RECT  6.740 -0.400 7.140 1.230 ;
        RECT  7.140 -0.400 7.150 1.030 ;
        RECT  7.150 -0.400 9.290 0.400 ;
        RECT  9.290 -0.400 9.300 1.200 ;
        RECT  9.300 -0.400 9.700 1.400 ;
        RECT  9.700 -0.400 9.710 1.200 ;
        RECT  9.710 -0.400 11.740 0.400 ;
        RECT  11.740 -0.400 11.750 0.670 ;
        RECT  11.750 -0.400 12.150 0.870 ;
        RECT  12.150 -0.400 12.160 0.670 ;
        RECT  12.160 -0.400 13.830 0.400 ;
        RECT  13.830 -0.400 14.230 0.560 ;
        RECT  14.230 -0.400 14.520 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.910 1.430 13.150 2.830 ;
        RECT  12.570 1.430 12.910 1.670 ;
        RECT  11.710 2.590 12.910 2.830 ;
        RECT  12.400 3.940 12.800 4.360 ;
        RECT  12.250 2.000 12.440 2.240 ;
        RECT  11.690 3.940 12.400 4.180 ;
        RECT  12.010 1.600 12.250 2.240 ;
        RECT  11.020 1.600 12.010 1.840 ;
        RECT  11.690 2.130 11.710 2.830 ;
        RECT  11.450 2.130 11.690 4.180 ;
        RECT  11.310 2.130 11.450 2.530 ;
        RECT  10.240 0.760 11.250 1.000 ;
        RECT  10.920 1.360 11.020 4.100 ;
        RECT  10.780 1.280 10.920 4.100 ;
        RECT  10.670 1.280 10.780 1.840 ;
        RECT  10.410 3.700 10.780 4.100 ;
        RECT  10.520 1.280 10.670 1.680 ;
        RECT  10.240 2.480 10.470 2.880 ;
        RECT  10.130 0.760 10.240 2.880 ;
        RECT  10.000 0.760 10.130 4.180 ;
        RECT  9.890 1.800 10.000 4.180 ;
        RECT  8.820 1.800 9.890 2.040 ;
        RECT  8.850 3.940 9.890 4.180 ;
        RECT  9.370 2.320 9.610 3.660 ;
        RECT  8.330 3.420 9.370 3.660 ;
        RECT  8.610 3.940 8.850 4.370 ;
        RECT  8.660 1.280 8.820 2.040 ;
        RECT  8.420 1.280 8.660 3.140 ;
        RECT  6.760 4.130 8.610 4.370 ;
        RECT  8.260 2.740 8.420 3.140 ;
        RECT  8.090 3.420 8.330 3.850 ;
        RECT  7.500 3.610 8.090 3.850 ;
        RECT  7.860 0.980 8.020 1.380 ;
        RECT  7.620 0.980 7.860 2.390 ;
        RECT  7.500 2.150 7.620 2.390 ;
        RECT  7.240 2.150 7.500 3.850 ;
        RECT  6.510 1.510 7.340 1.750 ;
        RECT  6.860 2.150 7.240 2.550 ;
        RECT  6.580 2.830 6.760 4.370 ;
        RECT  6.520 2.350 6.580 4.370 ;
        RECT  6.340 2.350 6.520 3.070 ;
        RECT  6.140 3.910 6.520 4.370 ;
        RECT  6.270 1.500 6.510 1.750 ;
        RECT  5.560 2.350 6.340 2.590 ;
        RECT  5.800 1.500 6.270 1.740 ;
        RECT  5.870 3.350 6.220 3.590 ;
        RECT  5.630 2.870 5.870 3.590 ;
        RECT  5.400 0.990 5.800 1.740 ;
        RECT  5.240 3.910 5.640 4.310 ;
        RECT  5.040 2.870 5.630 3.110 ;
        RECT  5.320 2.020 5.560 2.590 ;
        RECT  5.040 1.500 5.400 1.740 ;
        RECT  4.520 3.380 5.340 3.620 ;
        RECT  2.650 3.910 5.240 4.150 ;
        RECT  4.800 1.500 5.040 3.110 ;
        RECT  4.520 0.830 4.920 1.230 ;
        RECT  1.980 0.860 4.520 1.100 ;
        RECT  4.280 3.350 4.520 3.620 ;
        RECT  2.410 3.350 4.280 3.590 ;
        RECT  2.410 3.910 2.650 4.360 ;
        RECT  1.630 4.120 2.410 4.360 ;
        RECT  1.890 2.960 2.130 3.840 ;
        RECT  1.830 1.470 2.070 1.870 ;
        RECT  1.580 0.670 1.980 1.100 ;
        RECT  1.720 2.960 1.890 3.200 ;
        RECT  1.720 1.630 1.830 1.870 ;
        RECT  1.480 1.630 1.720 3.200 ;
        RECT  1.390 3.560 1.630 4.360 ;
        RECT  0.570 3.560 1.390 3.800 ;
        RECT  0.450 1.310 0.570 1.710 ;
        RECT  0.450 3.000 0.570 3.800 ;
        RECT  0.330 1.310 0.450 3.800 ;
        RECT  0.210 1.310 0.330 3.400 ;
        RECT  0.170 1.310 0.210 1.710 ;
        RECT  0.170 3.000 0.210 3.400 ;
    END
END SDFFNX1

MACRO SDFFHQXL
    CLASS CORE ;
    FOREIGN SDFFHQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.790 2.330 3.390 2.730 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.350 2.100 1.490 2.500 ;
        RECT  1.490 2.100 1.520 2.640 ;
        RECT  1.520 2.100 1.750 2.650 ;
        RECT  1.750 2.390 1.780 2.650 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.020 3.270 12.080 3.510 ;
        RECT  12.080 3.270 12.340 3.770 ;
        RECT  12.340 3.270 12.800 3.510 ;
        RECT  12.200 0.670 12.800 0.910 ;
        RECT  12.800 0.670 13.040 3.510 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.650 1.690 3.920 1.930 ;
        RECT  3.920 1.690 4.170 2.100 ;
        RECT  4.170 1.820 4.420 2.100 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.710 2.530 0.770 2.930 ;
        RECT  0.770 2.530 0.780 3.190 ;
        RECT  0.780 2.530 0.860 3.200 ;
        RECT  0.860 2.530 0.950 3.210 ;
        RECT  0.950 2.690 1.010 3.210 ;
        RECT  1.010 2.950 1.120 3.210 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.300 5.440 ;
        RECT  0.300 4.480 0.700 5.440 ;
        RECT  0.700 4.640 3.710 5.440 ;
        RECT  3.710 4.110 3.950 5.440 ;
        RECT  3.950 4.640 6.790 5.440 ;
        RECT  6.790 4.390 6.800 5.440 ;
        RECT  6.800 4.270 7.200 5.440 ;
        RECT  7.200 4.390 7.210 5.440 ;
        RECT  7.210 4.640 9.090 5.440 ;
        RECT  9.090 4.480 9.490 5.440 ;
        RECT  9.490 4.640 10.770 5.440 ;
        RECT  10.770 4.480 11.170 5.440 ;
        RECT  11.170 4.640 13.200 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.760 0.400 ;
        RECT  0.760 -0.400 1.120 1.730 ;
        RECT  1.120 1.370 1.460 1.730 ;
        RECT  1.120 -0.400 2.720 0.400 ;
        RECT  2.720 -0.400 3.120 0.560 ;
        RECT  3.120 -0.400 5.940 0.400 ;
        RECT  5.940 -0.400 5.950 0.730 ;
        RECT  5.950 -0.400 6.350 0.930 ;
        RECT  6.350 -0.400 6.360 0.730 ;
        RECT  6.360 -0.400 8.300 0.400 ;
        RECT  8.300 -0.400 8.310 0.750 ;
        RECT  8.310 -0.400 8.710 0.950 ;
        RECT  8.710 -0.400 8.720 0.750 ;
        RECT  8.720 -0.400 11.280 0.400 ;
        RECT  11.280 -0.400 11.290 0.670 ;
        RECT  11.290 -0.400 11.690 0.870 ;
        RECT  11.690 -0.400 11.700 0.670 ;
        RECT  11.700 -0.400 13.200 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.280 1.330 12.520 2.970 ;
        RECT  11.690 4.130 12.420 4.370 ;
        RECT  11.270 2.730 12.280 2.970 ;
        RECT  11.760 1.350 12.000 2.450 ;
        RECT  10.750 1.350 11.760 1.590 ;
        RECT  11.450 3.940 11.690 4.370 ;
        RECT  11.270 3.940 11.450 4.180 ;
        RECT  11.030 2.110 11.270 4.180 ;
        RECT  10.000 0.670 10.870 0.910 ;
        RECT  10.520 1.350 10.750 3.860 ;
        RECT  10.510 1.190 10.520 3.860 ;
        RECT  10.280 1.190 10.510 1.590 ;
        RECT  10.000 2.000 10.230 4.260 ;
        RECT  9.990 0.670 10.000 4.260 ;
        RECT  9.760 0.670 9.990 2.240 ;
        RECT  9.790 3.940 9.990 4.260 ;
        RECT  8.790 3.940 9.790 4.180 ;
        RECT  9.480 2.520 9.700 3.190 ;
        RECT  9.460 1.170 9.480 3.190 ;
        RECT  9.240 1.170 9.460 2.760 ;
        RECT  9.210 1.170 9.240 1.570 ;
        RECT  8.720 1.850 8.960 3.470 ;
        RECT  8.550 3.940 8.790 4.370 ;
        RECT  8.240 3.230 8.720 3.470 ;
        RECT  7.720 4.130 8.550 4.370 ;
        RECT  8.000 3.230 8.240 3.840 ;
        RECT  7.810 2.680 8.020 2.920 ;
        RECT  7.230 3.230 8.000 3.470 ;
        RECT  7.840 1.190 7.970 1.590 ;
        RECT  7.830 0.880 7.840 1.590 ;
        RECT  7.810 0.670 7.830 1.590 ;
        RECT  7.570 0.670 7.810 2.920 ;
        RECT  7.480 3.750 7.720 4.370 ;
        RECT  7.430 0.670 7.570 0.910 ;
        RECT  6.520 3.750 7.480 3.990 ;
        RECT  6.990 1.250 7.230 3.470 ;
        RECT  6.830 1.250 6.990 1.490 ;
        RECT  6.860 2.630 6.990 3.470 ;
        RECT  6.570 2.630 6.860 2.870 ;
        RECT  6.030 1.830 6.710 2.070 ;
        RECT  6.330 2.470 6.570 2.870 ;
        RECT  6.280 3.750 6.520 4.350 ;
        RECT  5.510 4.110 6.280 4.350 ;
        RECT  5.790 1.830 6.030 3.470 ;
        RECT  5.550 1.830 5.790 2.070 ;
        RECT  5.310 0.680 5.550 2.070 ;
        RECT  5.270 2.460 5.510 4.350 ;
        RECT  4.840 0.680 5.310 0.920 ;
        RECT  5.030 2.460 5.270 2.700 ;
        RECT  4.470 4.110 5.270 4.350 ;
        RECT  4.790 1.240 5.030 2.700 ;
        RECT  4.750 3.070 4.990 3.830 ;
        RECT  4.450 1.240 4.790 1.480 ;
        RECT  2.910 3.070 4.750 3.310 ;
        RECT  4.230 3.590 4.470 4.350 ;
        RECT  4.170 0.680 4.350 0.920 ;
        RECT  3.430 3.590 4.230 3.830 ;
        RECT  3.930 0.680 4.170 1.100 ;
        RECT  1.790 0.860 3.930 1.100 ;
        RECT  3.190 3.590 3.430 4.280 ;
        RECT  2.390 1.690 3.330 1.930 ;
        RECT  1.470 4.040 3.190 4.280 ;
        RECT  2.670 3.070 2.910 3.700 ;
        RECT  2.410 3.460 2.670 3.700 ;
        RECT  2.250 1.690 2.390 3.180 ;
        RECT  2.150 1.470 2.250 3.180 ;
        RECT  2.010 1.470 2.150 1.930 ;
        RECT  1.990 2.940 2.150 3.180 ;
        RECT  1.750 2.940 1.990 3.760 ;
        RECT  1.390 0.670 1.790 1.100 ;
        RECT  1.230 3.550 1.470 4.280 ;
        RECT  0.490 3.550 1.230 3.790 ;
        RECT  0.400 1.390 0.490 1.790 ;
        RECT  0.400 3.290 0.490 3.790 ;
        RECT  0.160 1.390 0.400 3.790 ;
    END
END SDFFHQXL

MACRO SDFFHQX4
    CLASS CORE ;
    FOREIGN SDFFHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFHQXL ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.020 2.740 3.420 3.140 ;
        RECT  3.420 2.740 4.070 2.980 ;
        RECT  4.070 2.420 4.160 2.980 ;
        RECT  4.160 2.390 4.310 2.980 ;
        RECT  4.310 2.390 4.410 2.660 ;
        RECT  4.410 2.390 4.420 2.650 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 2.390 2.280 2.650 ;
        RECT  2.280 2.010 2.440 2.650 ;
        RECT  2.440 2.010 2.520 2.640 ;
        RECT  2.520 2.010 3.800 2.420 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.010 2.730 17.270 3.740 ;
        RECT  16.990 0.660 17.270 1.640 ;
        RECT  17.270 0.660 17.390 3.740 ;
        RECT  17.390 1.400 17.410 3.740 ;
        RECT  17.410 1.400 17.510 3.220 ;
        RECT  17.510 1.820 17.710 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.390 1.370 4.730 1.630 ;
        RECT  4.730 1.270 5.080 1.630 ;
        RECT  5.080 1.280 5.160 1.630 ;
        RECT  5.160 1.370 5.170 1.630 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.690 1.970 0.860 2.370 ;
        RECT  0.860 1.830 1.110 2.370 ;
        RECT  1.110 1.830 1.120 2.090 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.030 5.440 ;
        RECT  1.030 4.370 1.040 5.440 ;
        RECT  1.040 4.250 1.440 5.440 ;
        RECT  1.440 4.370 1.450 5.440 ;
        RECT  1.450 4.640 3.920 5.440 ;
        RECT  3.920 4.480 4.320 5.440 ;
        RECT  4.320 4.640 6.830 5.440 ;
        RECT  6.830 4.480 7.230 5.440 ;
        RECT  7.230 4.640 9.170 5.440 ;
        RECT  9.170 3.910 9.180 5.440 ;
        RECT  9.180 3.710 9.580 5.440 ;
        RECT  9.580 3.910 9.590 5.440 ;
        RECT  9.590 4.640 12.940 5.440 ;
        RECT  12.940 3.980 12.950 5.440 ;
        RECT  12.950 3.860 13.350 5.440 ;
        RECT  13.350 3.980 13.360 5.440 ;
        RECT  13.360 4.640 14.720 5.440 ;
        RECT  14.720 4.480 15.120 5.440 ;
        RECT  15.120 4.640 16.430 5.440 ;
        RECT  16.250 3.300 16.430 3.700 ;
        RECT  16.430 3.300 16.670 5.440 ;
        RECT  16.670 4.640 17.830 5.440 ;
        RECT  17.830 3.820 18.230 5.440 ;
        RECT  18.230 4.640 18.480 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.030 0.400 ;
        RECT  1.030 -0.400 1.040 0.730 ;
        RECT  1.040 -0.400 1.440 0.930 ;
        RECT  1.440 -0.400 1.450 0.730 ;
        RECT  1.450 -0.400 3.340 0.400 ;
        RECT  3.340 -0.400 3.740 0.560 ;
        RECT  3.740 -0.400 6.690 0.400 ;
        RECT  6.690 -0.400 6.700 0.750 ;
        RECT  6.700 -0.400 7.100 0.950 ;
        RECT  7.100 -0.400 7.110 0.750 ;
        RECT  7.110 -0.400 9.190 0.400 ;
        RECT  9.190 -0.400 9.200 1.080 ;
        RECT  9.200 -0.400 9.600 1.200 ;
        RECT  9.600 -0.400 9.610 1.080 ;
        RECT  9.610 -0.400 13.050 0.400 ;
        RECT  13.050 -0.400 13.450 0.560 ;
        RECT  13.450 -0.400 14.600 0.400 ;
        RECT  14.600 -0.400 15.000 0.560 ;
        RECT  15.000 -0.400 16.220 0.400 ;
        RECT  16.220 -0.400 16.230 0.980 ;
        RECT  16.230 -0.400 16.630 1.470 ;
        RECT  16.630 -0.400 16.640 0.980 ;
        RECT  16.640 -0.400 17.800 0.400 ;
        RECT  17.800 -0.400 17.810 1.020 ;
        RECT  17.810 -0.400 18.210 1.220 ;
        RECT  18.210 -0.400 18.220 1.020 ;
        RECT  18.220 -0.400 18.230 0.560 ;
        RECT  18.230 -0.400 18.480 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  15.950 4.130 16.150 4.370 ;
        RECT  15.710 1.150 15.950 4.370 ;
        RECT  15.470 1.150 15.710 1.390 ;
        RECT  15.030 2.470 15.710 2.870 ;
        RECT  15.210 1.630 15.430 2.030 ;
        RECT  14.790 1.630 15.210 2.040 ;
        RECT  14.550 1.190 14.790 3.070 ;
        RECT  13.870 1.190 14.550 1.430 ;
        RECT  14.230 2.830 14.550 3.070 ;
        RECT  14.030 1.710 14.270 2.550 ;
        RECT  12.200 1.710 14.030 1.950 ;
        RECT  13.470 1.140 13.870 1.430 ;
        RECT  11.520 1.190 13.470 1.430 ;
        RECT  12.900 2.260 13.060 2.500 ;
        RECT  12.670 2.260 12.900 3.580 ;
        RECT  12.660 2.260 12.670 4.120 ;
        RECT  12.430 3.340 12.660 4.120 ;
        RECT  11.000 0.670 12.590 0.910 ;
        RECT  10.100 3.880 12.430 4.120 ;
        RECT  12.140 2.660 12.360 3.060 ;
        RECT  11.800 1.710 12.200 2.030 ;
        RECT  11.900 2.660 12.140 3.600 ;
        RECT  11.000 3.360 11.900 3.600 ;
        RECT  11.280 1.190 11.520 3.080 ;
        RECT  10.760 0.670 11.000 3.600 ;
        RECT  9.960 0.670 10.760 0.910 ;
        RECT  10.440 2.690 10.760 3.090 ;
        RECT  10.240 1.480 10.480 2.130 ;
        RECT  8.710 1.480 10.240 1.720 ;
        RECT  9.860 3.190 10.100 4.120 ;
        RECT  9.660 3.190 9.860 3.430 ;
        RECT  9.420 2.000 9.660 3.430 ;
        RECT  8.030 3.190 9.420 3.430 ;
        RECT  6.540 3.710 8.900 3.950 ;
        RECT  8.550 2.670 8.780 2.910 ;
        RECT  8.550 1.190 8.710 1.720 ;
        RECT  8.310 0.680 8.550 2.910 ;
        RECT  7.850 0.680 8.310 0.920 ;
        RECT  7.790 1.270 8.030 3.430 ;
        RECT  7.520 1.270 7.790 1.510 ;
        RECT  6.810 3.190 7.790 3.430 ;
        RECT  7.090 1.840 7.490 2.100 ;
        RECT  6.020 1.840 7.090 2.080 ;
        RECT  6.570 2.400 6.810 3.430 ;
        RECT  6.340 2.400 6.570 2.640 ;
        RECT  6.300 3.710 6.540 4.160 ;
        RECT  5.500 3.920 6.300 4.160 ;
        RECT  5.780 1.040 6.020 3.610 ;
        RECT  5.580 1.040 5.780 1.440 ;
        RECT  5.260 2.160 5.500 4.160 ;
        RECT  5.080 2.160 5.260 2.560 ;
        RECT  3.120 3.420 5.260 3.660 ;
        RECT  4.450 0.760 5.100 1.000 ;
        RECT  4.740 3.940 4.980 4.340 ;
        RECT  3.640 3.940 4.740 4.180 ;
        RECT  4.210 0.760 4.450 1.100 ;
        RECT  2.380 0.860 4.210 1.100 ;
        RECT  2.030 1.380 4.060 1.620 ;
        RECT  3.400 3.940 3.640 4.370 ;
        RECT  1.950 4.130 3.400 4.370 ;
        RECT  2.880 3.420 3.120 3.850 ;
        RECT  0.600 3.610 2.880 3.850 ;
        RECT  1.770 3.090 2.600 3.330 ;
        RECT  1.980 0.670 2.380 1.100 ;
        RECT  1.770 1.380 2.030 1.650 ;
        RECT  1.530 1.380 1.770 3.330 ;
        RECT  0.410 0.930 0.600 1.330 ;
        RECT  0.410 3.300 0.600 4.320 ;
        RECT  0.200 0.930 0.410 4.320 ;
        RECT  0.170 0.930 0.200 4.310 ;
    END
END SDFFHQX4

MACRO SDFFHQX2
    CLASS CORE ;
    FOREIGN SDFFHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFHQXL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.750 2.230 3.190 2.660 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.330 2.000 1.490 2.400 ;
        RECT  1.490 2.000 1.520 2.640 ;
        RECT  1.520 2.000 1.730 2.650 ;
        RECT  1.730 2.390 1.780 2.650 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.640 2.920 13.880 3.320 ;
        RECT  13.880 2.920 13.980 3.220 ;
        RECT  13.980 1.280 14.060 3.220 ;
        RECT  14.060 1.270 14.070 3.220 ;
        RECT  14.070 1.270 14.220 3.160 ;
        RECT  14.220 1.270 14.320 1.530 ;
        RECT  14.320 1.270 14.380 1.510 ;
        RECT  14.380 0.930 14.780 1.510 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.640 1.550 3.810 1.790 ;
        RECT  3.810 1.550 4.050 2.060 ;
        RECT  4.050 1.820 4.160 2.060 ;
        RECT  4.160 1.820 4.410 2.090 ;
        RECT  4.410 1.830 4.420 2.090 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.400 0.730 2.800 ;
        RECT  0.730 2.400 0.860 3.190 ;
        RECT  0.860 2.400 0.920 3.210 ;
        RECT  0.920 2.560 0.970 3.210 ;
        RECT  0.970 2.950 1.120 3.210 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.280 5.440 ;
        RECT  0.280 4.480 0.680 5.440 ;
        RECT  0.680 4.640 3.710 5.440 ;
        RECT  3.710 4.050 3.950 5.440 ;
        RECT  3.950 4.640 6.680 5.440 ;
        RECT  6.680 4.390 6.690 5.440 ;
        RECT  6.690 4.270 7.090 5.440 ;
        RECT  7.090 4.390 7.100 5.440 ;
        RECT  7.100 4.640 8.750 5.440 ;
        RECT  8.750 4.160 9.150 5.440 ;
        RECT  9.150 4.640 12.600 5.440 ;
        RECT  12.600 3.240 12.840 5.440 ;
        RECT  12.840 4.640 14.370 5.440 ;
        RECT  14.370 3.790 14.380 5.440 ;
        RECT  14.380 3.590 14.780 5.440 ;
        RECT  14.780 3.790 14.790 5.440 ;
        RECT  14.790 4.640 15.180 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.760 0.400 ;
        RECT  0.760 -0.400 1.120 1.730 ;
        RECT  1.120 1.370 1.340 1.730 ;
        RECT  1.120 -0.400 2.720 0.400 ;
        RECT  2.720 -0.400 3.120 0.560 ;
        RECT  3.120 -0.400 5.940 0.400 ;
        RECT  5.940 -0.400 5.950 0.730 ;
        RECT  5.950 -0.400 6.350 0.930 ;
        RECT  6.350 -0.400 6.360 0.730 ;
        RECT  6.360 -0.400 8.450 0.400 ;
        RECT  8.450 -0.400 8.850 0.560 ;
        RECT  8.850 -0.400 12.240 0.400 ;
        RECT  12.240 -0.400 12.640 0.560 ;
        RECT  12.640 -0.400 13.550 0.400 ;
        RECT  13.550 -0.400 13.950 0.560 ;
        RECT  13.950 -0.400 15.180 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  13.400 3.850 13.800 4.250 ;
        RECT  13.360 1.130 13.430 2.640 ;
        RECT  13.360 3.850 13.400 4.090 ;
        RECT  13.190 1.130 13.360 4.090 ;
        RECT  13.120 2.400 13.190 4.090 ;
        RECT  12.040 2.400 13.120 2.640 ;
        RECT  12.670 1.230 12.910 2.120 ;
        RECT  11.430 1.230 12.670 1.470 ;
        RECT  9.670 4.110 12.320 4.350 ;
        RECT  11.800 2.090 12.040 2.640 ;
        RECT  11.710 3.300 11.950 3.830 ;
        RECT  9.370 0.670 11.810 0.910 ;
        RECT  10.190 3.590 11.710 3.830 ;
        RECT  11.190 1.190 11.430 3.280 ;
        RECT  10.630 3.040 11.190 3.280 ;
        RECT  10.670 1.190 10.910 2.700 ;
        RECT  9.650 1.190 10.670 1.430 ;
        RECT  10.190 2.460 10.670 2.700 ;
        RECT  10.150 1.710 10.390 2.160 ;
        RECT  9.950 2.460 10.190 3.830 ;
        RECT  9.110 1.710 10.150 1.950 ;
        RECT  9.430 2.320 9.670 4.350 ;
        RECT  8.130 3.610 9.430 3.850 ;
        RECT  9.130 0.670 9.370 1.110 ;
        RECT  8.590 0.870 9.130 1.110 ;
        RECT  8.870 1.710 9.110 2.920 ;
        RECT  8.650 2.680 8.870 2.920 ;
        RECT  8.410 2.680 8.650 3.080 ;
        RECT  8.350 0.870 8.590 2.290 ;
        RECT  7.610 4.130 8.440 4.370 ;
        RECT  7.750 2.680 8.410 2.920 ;
        RECT  7.890 3.230 8.130 3.850 ;
        RECT  7.750 1.170 8.070 1.590 ;
        RECT  7.230 3.230 7.890 3.470 ;
        RECT  7.510 0.670 7.750 2.920 ;
        RECT  7.370 3.750 7.610 4.370 ;
        RECT  6.940 0.670 7.510 0.910 ;
        RECT  6.410 3.750 7.370 3.990 ;
        RECT  6.990 1.260 7.230 3.470 ;
        RECT  6.830 1.260 6.990 1.500 ;
        RECT  6.540 2.460 6.990 2.870 ;
        RECT  6.030 1.830 6.710 2.070 ;
        RECT  6.330 2.470 6.540 2.870 ;
        RECT  6.170 3.750 6.410 4.350 ;
        RECT  5.510 3.990 6.170 4.350 ;
        RECT  5.790 1.830 6.030 3.510 ;
        RECT  5.550 1.830 5.790 2.070 ;
        RECT  5.310 0.750 5.550 2.070 ;
        RECT  5.270 2.460 5.510 4.350 ;
        RECT  4.830 0.750 5.310 0.990 ;
        RECT  5.030 2.460 5.270 2.700 ;
        RECT  4.470 4.110 5.270 4.350 ;
        RECT  4.790 1.310 5.030 2.700 ;
        RECT  4.750 2.990 4.990 3.810 ;
        RECT  4.450 1.310 4.790 1.550 ;
        RECT  2.910 2.990 4.750 3.230 ;
        RECT  4.230 3.510 4.470 4.350 ;
        RECT  4.170 0.740 4.350 0.980 ;
        RECT  3.430 3.510 4.230 3.750 ;
        RECT  3.930 0.740 4.170 1.100 ;
        RECT  1.790 0.860 3.930 1.100 ;
        RECT  3.190 3.510 3.430 4.210 ;
        RECT  2.380 1.550 3.330 1.790 ;
        RECT  1.450 3.970 3.190 4.210 ;
        RECT  2.670 2.990 2.910 3.650 ;
        RECT  2.410 3.410 2.670 3.650 ;
        RECT  2.380 2.670 2.390 3.170 ;
        RECT  2.250 1.550 2.380 3.170 ;
        RECT  2.140 1.470 2.250 3.170 ;
        RECT  2.010 1.470 2.140 1.870 ;
        RECT  1.970 2.930 2.140 3.170 ;
        RECT  1.730 2.930 1.970 3.650 ;
        RECT  1.390 0.670 1.790 1.100 ;
        RECT  1.210 3.550 1.450 4.210 ;
        RECT  0.490 3.550 1.210 3.790 ;
        RECT  0.400 1.360 0.490 1.760 ;
        RECT  0.400 3.180 0.490 3.790 ;
        RECT  0.160 1.360 0.400 3.790 ;
    END
END SDFFHQX2

MACRO SDFFHQX1
    CLASS CORE ;
    FOREIGN SDFFHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFHQXL ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.750 2.230 3.190 2.660 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.330 2.000 1.490 2.400 ;
        RECT  1.490 2.000 1.520 2.640 ;
        RECT  1.520 2.000 1.730 2.650 ;
        RECT  1.730 2.390 1.780 2.650 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.960 3.250 11.990 3.490 ;
        RECT  11.990 3.250 12.080 3.760 ;
        RECT  12.080 3.250 12.340 3.770 ;
        RECT  12.340 3.250 12.430 3.760 ;
        RECT  12.430 3.250 12.800 3.490 ;
        RECT  12.140 0.670 12.800 0.910 ;
        RECT  12.800 0.670 13.040 3.490 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.650 1.470 3.930 1.870 ;
        RECT  3.930 1.470 4.160 2.080 ;
        RECT  4.160 1.470 4.170 2.090 ;
        RECT  4.170 1.830 4.420 2.090 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.530 0.730 2.930 ;
        RECT  0.730 2.530 0.860 3.190 ;
        RECT  0.860 2.530 0.920 3.210 ;
        RECT  0.920 2.690 0.970 3.210 ;
        RECT  0.970 2.950 1.120 3.210 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.280 5.440 ;
        RECT  0.280 4.480 0.680 5.440 ;
        RECT  0.680 4.640 3.710 5.440 ;
        RECT  3.710 4.050 3.950 5.440 ;
        RECT  3.950 4.640 6.790 5.440 ;
        RECT  6.790 4.390 6.800 5.440 ;
        RECT  6.800 4.270 7.200 5.440 ;
        RECT  7.200 4.390 7.210 5.440 ;
        RECT  7.210 4.640 9.090 5.440 ;
        RECT  9.090 4.480 9.490 5.440 ;
        RECT  9.490 4.640 10.770 5.440 ;
        RECT  10.770 4.480 11.170 5.440 ;
        RECT  11.170 4.640 13.200 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.760 0.400 ;
        RECT  0.760 -0.400 1.120 1.730 ;
        RECT  1.120 1.370 1.460 1.730 ;
        RECT  1.120 -0.400 2.720 0.400 ;
        RECT  2.720 -0.400 3.120 0.560 ;
        RECT  3.120 -0.400 5.940 0.400 ;
        RECT  5.940 -0.400 5.950 0.730 ;
        RECT  5.950 -0.400 6.350 0.930 ;
        RECT  6.350 -0.400 6.360 0.730 ;
        RECT  6.360 -0.400 8.330 0.400 ;
        RECT  8.330 -0.400 8.340 0.750 ;
        RECT  8.340 -0.400 8.740 0.950 ;
        RECT  8.740 -0.400 8.750 0.750 ;
        RECT  8.750 -0.400 11.280 0.400 ;
        RECT  11.280 -0.400 11.290 0.670 ;
        RECT  11.290 -0.400 11.690 0.870 ;
        RECT  11.690 -0.400 11.700 0.670 ;
        RECT  11.700 -0.400 13.200 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.280 1.350 12.520 2.970 ;
        RECT  11.690 4.130 12.420 4.370 ;
        RECT  11.270 2.730 12.280 2.970 ;
        RECT  11.760 1.350 12.000 2.450 ;
        RECT  10.750 1.350 11.760 1.590 ;
        RECT  11.450 3.940 11.690 4.370 ;
        RECT  11.270 3.940 11.450 4.180 ;
        RECT  11.030 2.080 11.270 4.180 ;
        RECT  10.000 0.680 10.920 0.920 ;
        RECT  10.520 1.350 10.750 3.760 ;
        RECT  10.510 1.200 10.520 3.760 ;
        RECT  10.280 1.200 10.510 1.600 ;
        RECT  10.000 2.000 10.230 4.260 ;
        RECT  9.990 0.680 10.000 4.260 ;
        RECT  9.760 0.680 9.990 2.240 ;
        RECT  9.790 3.940 9.990 4.260 ;
        RECT  8.790 3.940 9.790 4.180 ;
        RECT  9.480 2.520 9.700 3.430 ;
        RECT  9.460 1.050 9.480 3.430 ;
        RECT  9.240 1.050 9.460 2.760 ;
        RECT  8.760 2.070 9.000 3.470 ;
        RECT  8.550 3.940 8.790 4.370 ;
        RECT  8.240 3.230 8.760 3.470 ;
        RECT  7.720 4.130 8.550 4.370 ;
        RECT  8.000 3.230 8.240 3.840 ;
        RECT  7.810 2.680 8.020 2.920 ;
        RECT  7.230 3.230 8.000 3.470 ;
        RECT  7.810 1.210 7.970 1.610 ;
        RECT  7.570 0.670 7.810 2.920 ;
        RECT  7.480 3.750 7.720 4.370 ;
        RECT  6.970 0.670 7.570 0.910 ;
        RECT  6.410 3.750 7.480 3.990 ;
        RECT  6.990 1.250 7.230 3.470 ;
        RECT  6.830 1.250 6.990 1.490 ;
        RECT  6.860 2.630 6.990 3.470 ;
        RECT  6.570 2.630 6.860 2.870 ;
        RECT  6.030 1.830 6.710 2.070 ;
        RECT  6.330 2.470 6.570 2.870 ;
        RECT  6.170 3.750 6.410 4.350 ;
        RECT  6.010 3.990 6.170 4.350 ;
        RECT  5.790 1.830 6.030 3.510 ;
        RECT  5.510 3.990 6.010 4.230 ;
        RECT  5.550 1.830 5.790 2.070 ;
        RECT  5.310 0.750 5.550 2.070 ;
        RECT  5.270 2.460 5.510 4.230 ;
        RECT  4.830 0.750 5.310 0.990 ;
        RECT  5.030 2.460 5.270 2.700 ;
        RECT  4.470 3.990 5.270 4.230 ;
        RECT  4.790 1.310 5.030 2.700 ;
        RECT  4.750 2.990 4.990 3.700 ;
        RECT  4.450 1.310 4.790 1.550 ;
        RECT  2.910 2.990 4.750 3.230 ;
        RECT  4.230 3.510 4.470 4.230 ;
        RECT  4.170 0.740 4.350 0.980 ;
        RECT  3.430 3.510 4.230 3.750 ;
        RECT  3.930 0.740 4.170 1.100 ;
        RECT  1.790 0.860 3.930 1.100 ;
        RECT  3.190 3.510 3.430 4.220 ;
        RECT  2.930 1.470 3.330 1.870 ;
        RECT  1.450 3.980 3.190 4.220 ;
        RECT  2.380 1.550 2.930 1.790 ;
        RECT  2.670 2.990 2.910 3.690 ;
        RECT  2.410 3.450 2.670 3.690 ;
        RECT  2.380 2.670 2.390 3.170 ;
        RECT  2.250 1.550 2.380 3.170 ;
        RECT  2.140 1.470 2.250 3.170 ;
        RECT  2.010 1.470 2.140 1.870 ;
        RECT  1.970 2.930 2.140 3.170 ;
        RECT  1.730 2.930 1.970 3.650 ;
        RECT  1.390 0.670 1.790 1.100 ;
        RECT  1.210 3.550 1.450 4.220 ;
        RECT  0.490 3.550 1.210 3.790 ;
        RECT  0.400 1.360 0.490 1.790 ;
        RECT  0.400 3.390 0.490 3.790 ;
        RECT  0.160 1.360 0.400 3.790 ;
    END
END SDFFHQX1

MACRO SDFFXL
    CLASS CORE ;
    FOREIGN SDFFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.520 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.360 1.820 2.370 2.100 ;
        RECT  2.370 1.590 2.610 2.100 ;
        RECT  2.610 1.820 3.580 2.100 ;
        RECT  3.580 1.820 3.820 2.410 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.030 2.380 2.610 2.680 ;
        RECT  2.610 2.380 2.850 3.050 ;
        RECT  2.850 2.640 3.190 3.050 ;
        RECT  3.190 2.810 4.410 3.050 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.970 1.780 13.980 3.250 ;
        RECT  13.980 1.390 14.310 3.250 ;
        RECT  14.310 1.780 14.320 3.250 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.390 2.920 12.790 3.320 ;
        RECT  12.790 2.920 13.000 3.210 ;
        RECT  12.780 0.730 13.180 1.100 ;
        RECT  13.000 2.920 13.460 3.170 ;
        RECT  13.180 0.860 13.460 1.100 ;
        RECT  13.460 0.860 13.700 3.170 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.080 1.500 4.160 2.080 ;
        RECT  4.160 1.500 4.420 2.090 ;
        RECT  4.420 1.500 4.540 2.080 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.730 2.170 0.860 2.640 ;
        RECT  0.860 2.170 1.120 2.650 ;
        RECT  1.120 2.170 1.200 2.640 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.750 5.440 ;
        RECT  0.750 4.480 1.150 5.440 ;
        RECT  1.150 4.640 3.710 5.440 ;
        RECT  3.710 4.480 4.110 5.440 ;
        RECT  4.110 4.640 9.130 5.440 ;
        RECT  9.130 4.480 9.530 5.440 ;
        RECT  9.530 4.640 11.570 5.440 ;
        RECT  11.570 4.480 11.970 5.440 ;
        RECT  11.970 4.640 13.190 5.440 ;
        RECT  13.190 4.480 13.590 5.440 ;
        RECT  13.590 4.640 14.520 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.850 0.400 ;
        RECT  0.850 -0.400 1.250 0.560 ;
        RECT  1.250 -0.400 2.970 0.400 ;
        RECT  2.970 -0.400 3.370 0.560 ;
        RECT  3.370 -0.400 6.710 0.400 ;
        RECT  6.710 -0.400 7.110 1.180 ;
        RECT  7.110 -0.400 9.300 0.400 ;
        RECT  9.300 -0.400 9.700 1.490 ;
        RECT  9.700 -0.400 11.900 0.400 ;
        RECT  11.900 -0.400 12.300 1.070 ;
        RECT  12.300 -0.400 13.730 0.400 ;
        RECT  13.730 -0.400 14.130 0.560 ;
        RECT  14.130 -0.400 14.520 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.940 1.450 13.180 2.640 ;
        RECT  12.780 1.450 12.940 1.690 ;
        RECT  11.730 2.400 12.940 2.640 ;
        RECT  12.450 3.790 12.850 4.190 ;
        RECT  12.260 1.870 12.540 2.110 ;
        RECT  11.730 3.790 12.450 4.030 ;
        RECT  12.020 1.610 12.260 2.110 ;
        RECT  11.020 1.610 12.020 1.850 ;
        RECT  11.490 2.310 11.730 4.030 ;
        RECT  11.330 2.310 11.490 2.710 ;
        RECT  10.240 0.760 11.250 1.000 ;
        RECT  10.780 1.290 11.020 4.220 ;
        RECT  10.520 1.290 10.780 1.690 ;
        RECT  10.470 3.820 10.780 4.220 ;
        RECT  10.240 2.610 10.480 3.010 ;
        RECT  10.190 0.760 10.240 3.010 ;
        RECT  10.000 0.760 10.190 4.180 ;
        RECT  8.950 1.800 10.000 2.040 ;
        RECT  9.950 2.770 10.000 4.180 ;
        RECT  8.850 3.940 9.950 4.180 ;
        RECT  9.430 2.320 9.670 3.660 ;
        RECT  8.330 3.420 9.430 3.660 ;
        RECT  8.710 1.800 8.950 2.460 ;
        RECT  8.610 3.940 8.850 4.370 ;
        RECT  8.680 1.260 8.820 1.500 ;
        RECT  8.460 2.770 8.730 3.170 ;
        RECT  8.460 0.670 8.680 1.500 ;
        RECT  6.760 4.130 8.610 4.370 ;
        RECT  8.330 0.670 8.460 3.170 ;
        RECT  8.220 0.670 8.330 3.090 ;
        RECT  8.090 3.420 8.330 3.840 ;
        RECT  7.500 3.600 8.090 3.840 ;
        RECT  7.670 1.000 7.910 2.390 ;
        RECT  7.500 2.150 7.670 2.390 ;
        RECT  7.240 2.150 7.500 3.840 ;
        RECT  5.770 1.500 7.390 1.740 ;
        RECT  6.860 2.150 7.240 2.550 ;
        RECT  6.580 2.890 6.760 4.370 ;
        RECT  6.520 2.350 6.580 4.370 ;
        RECT  6.340 2.350 6.520 3.130 ;
        RECT  6.110 3.910 6.520 4.370 ;
        RECT  5.570 2.350 6.340 2.590 ;
        RECT  5.900 3.410 6.200 3.650 ;
        RECT  2.710 3.910 6.110 4.150 ;
        RECT  5.660 2.870 5.900 3.650 ;
        RECT  5.370 0.860 5.770 1.740 ;
        RECT  5.050 2.870 5.660 3.110 ;
        RECT  5.330 2.020 5.570 2.590 ;
        RECT  2.470 3.370 5.380 3.610 ;
        RECT  5.050 1.500 5.370 1.740 ;
        RECT  4.810 1.500 5.050 3.110 ;
        RECT  4.490 0.820 4.890 1.220 ;
        RECT  1.980 0.860 4.490 1.100 ;
        RECT  2.470 3.910 2.710 4.360 ;
        RECT  1.670 4.120 2.470 4.360 ;
        RECT  1.950 2.950 2.190 3.840 ;
        RECT  1.800 1.460 2.040 1.870 ;
        RECT  1.580 0.660 1.980 1.100 ;
        RECT  1.760 2.950 1.950 3.190 ;
        RECT  1.760 1.630 1.800 1.870 ;
        RECT  1.520 1.630 1.760 3.190 ;
        RECT  1.430 3.540 1.670 4.360 ;
        RECT  0.570 3.540 1.430 3.780 ;
        RECT  0.410 1.320 0.570 1.720 ;
        RECT  0.410 2.930 0.570 3.780 ;
        RECT  0.330 1.320 0.410 3.780 ;
        RECT  0.170 1.320 0.330 3.330 ;
    END
END SDFFXL

MACRO SDFFX4
    CLASS CORE ;
    FOREIGN SDFFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFXL ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.950 2.870 3.210 ;
        RECT  2.870 2.710 2.880 3.210 ;
        RECT  2.880 2.540 3.100 3.210 ;
        RECT  3.100 2.540 3.280 3.200 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.990 2.220 2.360 2.660 ;
        RECT  2.360 2.020 2.610 2.660 ;
        RECT  2.610 2.020 3.560 2.260 ;
        RECT  3.560 2.020 3.800 2.840 ;
        RECT  3.800 2.600 3.940 2.840 ;
        RECT  3.940 2.600 4.340 3.000 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.930 1.820 18.100 3.220 ;
        RECT  18.100 1.410 18.110 3.220 ;
        RECT  18.110 1.210 18.310 3.220 ;
        RECT  18.310 1.210 18.510 3.270 ;
        RECT  18.510 1.410 18.520 3.270 ;
        RECT  18.520 2.870 18.710 3.270 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.610 1.820 16.760 3.220 ;
        RECT  16.760 1.410 16.770 3.220 ;
        RECT  16.770 1.210 17.170 3.270 ;
        RECT  17.170 1.410 17.180 3.070 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.070 1.510 4.510 2.100 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.710 1.920 0.860 2.640 ;
        RECT  0.860 1.920 1.120 2.650 ;
        RECT  1.120 1.920 1.180 2.640 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 4.480 1.390 5.440 ;
        RECT  1.390 4.640 6.930 5.440 ;
        RECT  6.930 4.480 7.330 5.440 ;
        RECT  7.330 4.640 9.480 5.440 ;
        RECT  9.480 4.480 9.880 5.440 ;
        RECT  9.880 4.640 11.980 5.440 ;
        RECT  11.980 4.140 12.380 5.440 ;
        RECT  12.380 4.640 14.530 5.440 ;
        RECT  14.530 4.480 14.930 5.440 ;
        RECT  14.930 4.640 16.130 5.440 ;
        RECT  16.130 4.070 16.530 5.440 ;
        RECT  16.530 4.640 17.510 5.440 ;
        RECT  17.510 4.070 17.910 5.440 ;
        RECT  17.910 4.640 18.950 5.440 ;
        RECT  18.950 4.070 19.350 5.440 ;
        RECT  19.350 4.640 19.800 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.930 0.400 ;
        RECT  0.930 -0.400 1.330 1.030 ;
        RECT  1.330 -0.400 3.010 0.400 ;
        RECT  3.010 -0.400 3.410 0.560 ;
        RECT  3.410 -0.400 6.680 0.400 ;
        RECT  6.680 -0.400 7.080 1.300 ;
        RECT  7.080 -0.400 9.530 0.400 ;
        RECT  9.530 -0.400 9.930 1.400 ;
        RECT  9.930 -0.400 11.970 0.400 ;
        RECT  11.970 -0.400 12.370 1.300 ;
        RECT  12.370 -0.400 14.560 0.400 ;
        RECT  14.560 -0.400 14.960 0.560 ;
        RECT  14.960 -0.400 16.130 0.400 ;
        RECT  16.130 -0.400 16.530 0.930 ;
        RECT  16.530 -0.400 17.440 0.400 ;
        RECT  17.440 -0.400 17.840 0.930 ;
        RECT  17.840 -0.400 18.750 0.400 ;
        RECT  18.750 -0.400 19.150 0.930 ;
        RECT  19.150 -0.400 19.800 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  18.990 2.190 19.230 3.790 ;
        RECT  18.820 2.190 18.990 2.590 ;
        RECT  16.340 3.550 18.990 3.790 ;
        RECT  16.100 1.260 16.340 3.790 ;
        RECT  15.780 1.260 16.100 1.500 ;
        RECT  15.260 3.390 16.100 3.790 ;
        RECT  15.580 2.260 15.820 3.050 ;
        RECT  15.380 1.100 15.780 1.500 ;
        RECT  14.410 2.810 15.580 3.050 ;
        RECT  14.930 1.260 15.380 1.500 ;
        RECT  14.690 1.260 14.930 2.520 ;
        RECT  14.170 0.980 14.410 3.860 ;
        RECT  12.930 0.980 14.170 1.220 ;
        RECT  13.640 3.620 14.170 3.860 ;
        RECT  13.600 1.510 13.840 2.910 ;
        RECT  13.240 3.620 13.640 4.020 ;
        RECT  13.400 2.670 13.600 2.910 ;
        RECT  12.990 2.670 13.400 3.340 ;
        RECT  11.160 3.620 13.240 3.860 ;
        RECT  10.970 3.100 12.990 3.340 ;
        RECT  12.690 0.980 12.930 1.830 ;
        RECT  11.150 1.590 12.690 1.830 ;
        RECT  11.730 2.110 12.130 2.510 ;
        RECT  10.180 2.110 11.730 2.350 ;
        RECT  10.760 3.620 11.160 4.110 ;
        RECT  10.750 1.240 11.150 1.830 ;
        RECT  10.560 2.640 10.970 3.340 ;
        RECT  10.480 3.100 10.560 3.340 ;
        RECT  10.240 3.100 10.480 4.180 ;
        RECT  9.470 3.940 10.240 4.180 ;
        RECT  10.100 1.920 10.180 2.630 ;
        RECT  9.770 1.680 10.100 2.630 ;
        RECT  9.250 1.680 9.770 1.920 ;
        RECT  9.230 2.210 9.470 4.180 ;
        RECT  9.010 0.760 9.250 1.920 ;
        RECT  9.030 2.210 9.230 2.610 ;
        RECT  6.550 3.940 9.230 4.180 ;
        RECT  7.840 0.760 9.010 1.000 ;
        RECT  8.730 3.030 8.950 3.430 ;
        RECT  8.490 1.280 8.730 3.430 ;
        RECT  8.330 1.280 8.490 2.260 ;
        RECT  8.130 1.860 8.330 2.260 ;
        RECT  7.840 3.420 8.150 3.660 ;
        RECT  7.600 0.760 7.840 3.660 ;
        RECT  7.440 1.100 7.600 1.500 ;
        RECT  7.190 2.660 7.600 2.900 ;
        RECT  6.920 1.830 7.320 2.180 ;
        RECT  6.790 2.580 7.190 2.980 ;
        RECT  6.070 1.830 6.920 2.070 ;
        RECT  6.510 3.940 6.550 4.240 ;
        RECT  6.270 2.350 6.510 4.240 ;
        RECT  5.530 2.350 6.270 2.590 ;
        RECT  4.330 4.000 6.270 4.240 ;
        RECT  5.830 1.420 6.070 2.070 ;
        RECT  5.750 2.880 5.990 3.690 ;
        RECT  5.710 1.420 5.830 1.660 ;
        RECT  5.020 2.880 5.750 3.120 ;
        RECT  5.310 0.690 5.710 1.660 ;
        RECT  5.290 1.940 5.530 2.590 ;
        RECT  5.020 1.420 5.310 1.660 ;
        RECT  3.800 3.400 5.310 3.640 ;
        RECT  4.780 1.420 5.020 3.120 ;
        RECT  4.430 0.720 4.830 1.120 ;
        RECT  3.930 0.880 4.430 1.120 ;
        RECT  4.090 4.000 4.330 4.300 ;
        RECT  1.910 4.060 4.090 4.300 ;
        RECT  3.690 0.880 3.930 1.220 ;
        RECT  2.070 1.500 3.800 1.740 ;
        RECT  3.560 3.400 3.800 3.770 ;
        RECT  2.070 0.980 3.690 1.220 ;
        RECT  2.470 3.530 3.560 3.770 ;
        RECT  1.910 2.940 2.480 3.180 ;
        RECT  1.670 0.760 2.070 1.220 ;
        RECT  1.720 1.500 2.070 1.900 ;
        RECT  1.720 2.940 1.910 3.260 ;
        RECT  1.670 3.840 1.910 4.300 ;
        RECT  1.480 1.500 1.720 3.260 ;
        RECT  0.570 3.840 1.670 4.080 ;
        RECT  0.430 1.200 0.570 1.600 ;
        RECT  0.430 3.110 0.570 4.090 ;
        RECT  0.190 1.200 0.430 4.090 ;
        RECT  0.170 1.200 0.190 1.600 ;
        RECT  0.170 3.110 0.190 4.090 ;
    END
END SDFFX4

MACRO SDFFX2
    CLASS CORE ;
    FOREIGN SDFFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.360 1.820 2.370 2.100 ;
        RECT  2.370 1.590 2.610 2.100 ;
        RECT  2.610 1.820 3.520 2.100 ;
        RECT  3.520 1.820 3.760 2.410 ;
        RECT  3.760 1.820 3.780 2.100 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.000 2.390 2.590 2.660 ;
        RECT  2.590 2.390 2.830 3.060 ;
        RECT  2.830 2.820 4.290 3.060 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.530 3.130 16.610 4.110 ;
        RECT  16.450 0.730 16.610 1.710 ;
        RECT  16.610 0.730 16.850 4.110 ;
        RECT  16.850 2.390 16.960 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.700 0.690 15.110 1.100 ;
        RECT  14.650 3.130 15.480 3.530 ;
        RECT  15.110 0.860 15.480 1.100 ;
        RECT  15.480 0.860 15.720 3.530 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 1.560 4.510 2.090 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.730 2.170 0.860 2.640 ;
        RECT  0.860 2.170 1.120 2.650 ;
        RECT  1.120 2.170 1.180 2.640 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.730 5.440 ;
        RECT  0.730 4.480 1.130 5.440 ;
        RECT  1.130 4.640 3.740 5.440 ;
        RECT  3.740 4.480 4.140 5.440 ;
        RECT  4.140 4.640 8.950 5.440 ;
        RECT  8.950 4.480 9.350 5.440 ;
        RECT  9.350 4.640 11.500 5.440 ;
        RECT  11.500 4.480 11.900 5.440 ;
        RECT  11.900 4.640 13.710 5.440 ;
        RECT  13.710 4.480 14.110 5.440 ;
        RECT  14.110 4.640 15.530 5.440 ;
        RECT  15.530 4.480 15.930 5.440 ;
        RECT  15.930 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.300 0.400 ;
        RECT  0.300 -0.400 0.700 0.560 ;
        RECT  0.700 -0.400 2.890 0.400 ;
        RECT  2.890 -0.400 3.290 0.560 ;
        RECT  3.290 -0.400 6.680 0.400 ;
        RECT  6.680 -0.400 7.080 1.250 ;
        RECT  7.080 -0.400 9.300 0.400 ;
        RECT  9.300 -0.400 9.700 1.390 ;
        RECT  9.700 -0.400 11.740 0.400 ;
        RECT  11.740 -0.400 12.140 1.390 ;
        RECT  12.140 -0.400 13.930 0.400 ;
        RECT  13.930 -0.400 14.330 0.990 ;
        RECT  14.330 -0.400 15.630 0.400 ;
        RECT  15.630 -0.400 16.030 0.560 ;
        RECT  16.030 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.000 2.170 16.240 4.090 ;
        RECT  15.050 3.850 16.000 4.090 ;
        RECT  14.980 1.380 15.070 1.780 ;
        RECT  14.650 3.850 15.050 4.320 ;
        RECT  14.740 1.380 14.980 2.800 ;
        RECT  14.370 2.560 14.740 2.800 ;
        RECT  14.370 3.850 14.650 4.090 ;
        RECT  14.250 1.600 14.490 2.320 ;
        RECT  14.130 2.560 14.370 4.090 ;
        RECT  13.250 1.600 14.250 1.840 ;
        RECT  13.770 2.560 14.130 2.850 ;
        RECT  13.530 2.180 13.770 2.850 ;
        RECT  13.010 1.600 13.250 3.640 ;
        RECT  12.990 1.600 13.010 1.920 ;
        RECT  12.640 3.400 13.010 3.640 ;
        RECT  12.590 1.110 12.990 1.920 ;
        RECT  12.490 2.410 12.730 2.860 ;
        RECT  12.240 3.400 12.640 3.800 ;
        RECT  10.920 1.680 12.590 1.920 ;
        RECT  10.380 2.620 12.490 2.860 ;
        RECT  10.620 3.520 12.240 3.760 ;
        RECT  10.680 1.240 10.920 1.920 ;
        RECT  10.520 1.240 10.680 1.640 ;
        RECT  10.220 3.520 10.620 3.920 ;
        RECT  10.240 2.620 10.380 3.240 ;
        RECT  10.000 1.680 10.240 3.240 ;
        RECT  8.770 1.680 10.000 1.920 ;
        RECT  9.970 2.620 10.000 3.240 ;
        RECT  9.610 3.000 9.970 3.240 ;
        RECT  9.240 2.320 9.640 2.720 ;
        RECT  9.370 3.000 9.610 4.180 ;
        RECT  8.660 3.940 9.370 4.180 ;
        RECT  9.080 2.480 9.240 2.720 ;
        RECT  8.840 2.480 9.080 3.660 ;
        RECT  8.140 3.420 8.840 3.660 ;
        RECT  8.420 1.070 8.820 1.310 ;
        RECT  8.420 3.940 8.660 4.370 ;
        RECT  8.420 2.740 8.560 3.140 ;
        RECT  8.180 1.070 8.420 3.140 ;
        RECT  6.730 4.130 8.420 4.370 ;
        RECT  8.130 2.020 8.180 3.140 ;
        RECT  7.740 3.420 8.140 3.800 ;
        RECT  7.740 0.910 7.900 1.310 ;
        RECT  7.500 0.910 7.740 3.800 ;
        RECT  6.640 2.290 7.500 2.530 ;
        RECT  6.820 1.500 7.220 1.810 ;
        RECT  5.710 1.500 6.820 1.740 ;
        RECT  6.490 2.880 6.730 4.370 ;
        RECT  6.360 2.880 6.490 3.120 ;
        RECT  6.100 3.920 6.490 4.370 ;
        RECT  6.120 2.350 6.360 3.120 ;
        RECT  5.840 3.390 6.200 3.630 ;
        RECT  5.540 2.350 6.120 2.590 ;
        RECT  2.740 3.920 6.100 4.160 ;
        RECT  5.600 2.870 5.840 3.630 ;
        RECT  5.310 1.050 5.710 1.740 ;
        RECT  5.020 2.870 5.600 3.110 ;
        RECT  5.300 2.020 5.540 2.590 ;
        RECT  2.410 3.390 5.320 3.630 ;
        RECT  5.020 1.500 5.310 1.740 ;
        RECT  4.780 1.500 5.020 3.110 ;
        RECT  4.430 0.830 4.830 1.230 ;
        RECT  1.950 0.860 4.430 1.100 ;
        RECT  2.500 3.920 2.740 4.320 ;
        RECT  1.640 4.080 2.500 4.320 ;
        RECT  1.900 2.950 2.140 3.840 ;
        RECT  1.770 1.460 2.010 1.870 ;
        RECT  1.550 0.660 1.950 1.100 ;
        RECT  1.720 2.950 1.900 3.190 ;
        RECT  1.720 1.630 1.770 1.870 ;
        RECT  1.480 1.630 1.720 3.190 ;
        RECT  1.400 3.870 1.640 4.320 ;
        RECT  0.570 3.870 1.400 4.110 ;
        RECT  0.450 1.320 0.570 1.720 ;
        RECT  0.450 3.000 0.570 4.110 ;
        RECT  0.330 1.320 0.450 4.110 ;
        RECT  0.210 1.320 0.330 3.400 ;
        RECT  0.170 1.320 0.210 1.720 ;
        RECT  0.170 3.000 0.210 3.400 ;
    END
END SDFFX2

MACRO SDFFX1
    CLASS CORE ;
    FOREIGN SDFFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ SDFFXL ;
    SIZE 14.520 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.330 1.820 2.340 2.100 ;
        RECT  2.340 1.590 2.580 2.100 ;
        RECT  2.580 1.820 3.520 2.100 ;
        RECT  3.520 1.820 3.760 2.410 ;
        RECT  3.760 1.820 3.780 2.100 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.030 2.380 2.590 2.680 ;
        RECT  2.590 2.380 2.830 3.050 ;
        RECT  2.830 2.810 4.290 3.050 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.820 3.570 14.020 3.810 ;
        RECT  14.020 1.540 14.030 3.810 ;
        RECT  14.030 1.320 14.310 3.810 ;
        RECT  14.310 2.390 14.320 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.260 3.050 12.650 3.450 ;
        RECT  12.650 3.050 12.740 3.740 ;
        RECT  12.510 0.690 12.910 1.100 ;
        RECT  12.740 3.050 13.000 3.770 ;
        RECT  13.000 3.050 13.090 3.740 ;
        RECT  13.090 3.050 13.460 3.290 ;
        RECT  12.910 0.860 13.460 1.100 ;
        RECT  13.460 0.860 13.700 3.290 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.080 1.500 4.160 2.080 ;
        RECT  4.160 1.500 4.420 2.090 ;
        RECT  4.420 1.500 4.510 2.080 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.730 2.170 0.860 2.640 ;
        RECT  0.860 2.170 1.120 2.650 ;
        RECT  1.120 2.170 1.200 2.640 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.730 5.440 ;
        RECT  0.730 4.480 1.130 5.440 ;
        RECT  1.130 4.640 3.750 5.440 ;
        RECT  3.750 4.480 4.150 5.440 ;
        RECT  4.150 4.640 9.130 5.440 ;
        RECT  9.130 4.480 9.530 5.440 ;
        RECT  9.530 4.640 11.440 5.440 ;
        RECT  11.440 4.480 11.840 5.440 ;
        RECT  11.840 4.640 13.060 5.440 ;
        RECT  13.060 4.480 13.460 5.440 ;
        RECT  13.460 4.640 14.520 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.300 0.400 ;
        RECT  0.300 -0.400 0.700 0.560 ;
        RECT  0.700 -0.400 2.890 0.400 ;
        RECT  2.890 -0.400 3.290 0.560 ;
        RECT  3.290 -0.400 6.680 0.400 ;
        RECT  6.680 -0.400 7.080 1.160 ;
        RECT  7.080 -0.400 9.300 0.400 ;
        RECT  9.300 -0.400 9.700 1.390 ;
        RECT  9.700 -0.400 11.750 0.400 ;
        RECT  11.750 -0.400 12.150 0.860 ;
        RECT  12.150 -0.400 13.800 0.400 ;
        RECT  13.800 -0.400 14.200 0.560 ;
        RECT  14.200 -0.400 14.520 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.940 1.420 13.180 2.770 ;
        RECT  12.570 1.420 12.940 1.660 ;
        RECT  11.710 2.530 12.940 2.770 ;
        RECT  12.380 4.050 12.660 4.290 ;
        RECT  12.250 2.000 12.410 2.240 ;
        RECT  12.140 3.940 12.380 4.290 ;
        RECT  12.010 1.600 12.250 2.240 ;
        RECT  11.690 3.940 12.140 4.180 ;
        RECT  10.920 1.600 12.010 1.840 ;
        RECT  11.690 2.130 11.710 2.770 ;
        RECT  11.450 2.130 11.690 4.180 ;
        RECT  11.310 2.130 11.450 2.530 ;
        RECT  10.240 0.760 11.250 1.000 ;
        RECT  10.910 1.290 10.920 1.840 ;
        RECT  10.670 1.290 10.910 4.370 ;
        RECT  10.520 1.290 10.670 1.690 ;
        RECT  10.410 3.970 10.670 4.370 ;
        RECT  10.240 2.310 10.280 2.710 ;
        RECT  10.170 0.760 10.240 2.710 ;
        RECT  10.000 0.760 10.170 4.230 ;
        RECT  8.770 1.640 10.000 1.880 ;
        RECT  9.930 2.390 10.000 4.230 ;
        RECT  8.850 3.990 9.930 4.230 ;
        RECT  9.320 2.240 9.560 3.750 ;
        RECT  8.330 3.510 9.320 3.750 ;
        RECT  8.610 3.990 8.850 4.370 ;
        RECT  8.420 0.850 8.820 1.250 ;
        RECT  6.710 4.130 8.610 4.370 ;
        RECT  8.380 2.800 8.560 3.200 ;
        RECT  8.380 1.010 8.420 1.250 ;
        RECT  8.140 1.010 8.380 3.200 ;
        RECT  8.090 3.510 8.330 3.850 ;
        RECT  7.480 3.610 8.090 3.850 ;
        RECT  7.640 0.760 7.880 2.270 ;
        RECT  7.480 2.030 7.640 2.270 ;
        RECT  7.210 2.030 7.480 3.850 ;
        RECT  5.710 1.500 7.340 1.740 ;
        RECT  6.810 2.150 7.210 2.550 ;
        RECT  6.490 2.890 6.710 4.370 ;
        RECT  6.470 2.350 6.490 4.370 ;
        RECT  6.250 2.350 6.470 3.130 ;
        RECT  6.120 3.920 6.470 4.370 ;
        RECT  5.530 2.350 6.250 2.590 ;
        RECT  5.840 3.400 6.200 3.640 ;
        RECT  2.730 3.920 6.120 4.160 ;
        RECT  5.600 2.870 5.840 3.640 ;
        RECT  5.310 0.990 5.710 1.740 ;
        RECT  5.020 2.870 5.600 3.110 ;
        RECT  5.290 2.020 5.530 2.590 ;
        RECT  2.410 3.380 5.320 3.620 ;
        RECT  5.020 1.500 5.310 1.740 ;
        RECT  4.780 1.500 5.020 3.110 ;
        RECT  4.670 0.970 4.830 1.210 ;
        RECT  4.430 0.860 4.670 1.210 ;
        RECT  2.610 0.860 4.430 1.100 ;
        RECT  2.490 3.920 2.730 4.320 ;
        RECT  2.370 0.670 2.610 1.100 ;
        RECT  1.630 4.080 2.490 4.320 ;
        RECT  1.550 0.670 2.370 0.910 ;
        RECT  1.890 2.950 2.130 3.840 ;
        RECT  1.790 1.460 2.010 1.860 ;
        RECT  1.790 2.950 1.890 3.190 ;
        RECT  1.550 1.460 1.790 3.190 ;
        RECT  1.390 3.900 1.630 4.320 ;
        RECT  0.570 3.900 1.390 4.140 ;
        RECT  0.450 1.310 0.570 1.710 ;
        RECT  0.450 3.000 0.570 4.140 ;
        RECT  0.330 1.310 0.450 4.140 ;
        RECT  0.210 1.310 0.330 3.400 ;
        RECT  0.170 1.310 0.210 1.710 ;
        RECT  0.170 3.000 0.210 3.400 ;
    END
END SDFFX1

MACRO RSLATNXL
    CLASS CORE ;
    FOREIGN RSLATNXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.070 2.370 3.230 2.610 ;
        RECT  3.230 1.850 3.470 2.610 ;
        RECT  3.470 1.850 3.500 2.090 ;
        RECT  3.500 1.830 3.760 2.090 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.910 2.370 4.510 2.670 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.140 2.950 6.150 3.210 ;
        RECT  6.150 2.870 6.810 3.270 ;
        RECT  6.690 1.390 6.810 1.790 ;
        RECT  6.810 2.640 6.850 3.270 ;
        RECT  6.810 1.390 6.850 1.840 ;
        RECT  6.850 1.390 7.090 3.270 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.160 3.510 0.170 4.130 ;
        RECT  0.170 1.390 0.410 4.130 ;
        RECT  0.410 1.390 0.450 1.840 ;
        RECT  0.450 1.390 0.570 1.790 ;
        RECT  0.410 3.510 0.580 4.130 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.980 5.440 ;
        RECT  0.980 3.900 0.990 5.440 ;
        RECT  0.990 3.700 1.390 5.440 ;
        RECT  1.390 3.900 1.400 5.440 ;
        RECT  1.400 4.640 2.780 5.440 ;
        RECT  2.780 4.480 3.760 5.440 ;
        RECT  3.760 4.640 6.080 5.440 ;
        RECT  6.080 4.480 6.480 5.440 ;
        RECT  6.480 4.640 7.260 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.280 0.400 ;
        RECT  0.280 -0.400 0.680 0.560 ;
        RECT  0.680 -0.400 2.650 0.400 ;
        RECT  2.650 -0.400 3.050 0.560 ;
        RECT  3.050 -0.400 4.290 0.400 ;
        RECT  4.290 -0.400 4.690 0.560 ;
        RECT  4.690 -0.400 6.580 0.400 ;
        RECT  6.580 -0.400 6.980 0.560 ;
        RECT  6.980 -0.400 7.260 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.250 2.090 6.570 2.490 ;
        RECT  6.010 0.800 6.250 2.490 ;
        RECT  5.610 0.800 6.010 1.040 ;
        RECT  5.760 2.250 6.010 2.490 ;
        RECT  5.520 2.250 5.760 3.850 ;
        RECT  4.930 1.330 5.740 1.570 ;
        RECT  5.210 0.760 5.610 1.040 ;
        RECT  5.210 3.610 5.520 3.850 ;
        RECT  5.020 2.430 5.210 2.830 ;
        RECT  4.810 3.610 5.210 4.010 ;
        RECT  4.780 1.850 5.020 3.190 ;
        RECT  4.690 0.860 4.930 1.570 ;
        RECT  2.490 3.770 4.810 4.010 ;
        RECT  4.410 1.850 4.780 2.090 ;
        RECT  4.290 2.950 4.780 3.190 ;
        RECT  2.070 0.860 4.690 1.100 ;
        RECT  4.170 1.380 4.410 2.090 ;
        RECT  2.790 2.940 3.850 3.180 ;
        RECT  2.790 1.380 2.870 1.790 ;
        RECT  2.630 1.380 2.790 3.180 ;
        RECT  2.550 1.550 2.630 3.180 ;
        RECT  1.370 1.550 2.550 1.950 ;
        RECT  2.100 3.770 2.490 4.300 ;
        RECT  2.090 3.900 2.100 4.300 ;
        RECT  1.670 0.790 2.070 1.190 ;
        RECT  1.510 2.910 1.910 3.310 ;
        RECT  1.090 0.950 1.670 1.190 ;
        RECT  1.090 2.910 1.510 3.150 ;
        RECT  0.850 0.950 1.090 3.150 ;
        RECT  0.730 2.070 0.850 2.470 ;
    END
END RSLATNXL

MACRO RSLATNX4
    CLASS CORE ;
    FOREIGN RSLATNX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ RSLATNXL ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.800 1.830 2.200 2.470 ;
        RECT  2.200 1.830 2.440 2.090 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  10.040 1.910 10.100 2.310 ;
        RECT  10.100 1.830 10.360 2.310 ;
        RECT  10.360 1.910 10.440 2.310 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.170 1.270 11.330 3.150 ;
        RECT  11.330 1.260 11.570 3.150 ;
        RECT  11.570 1.260 11.770 2.660 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.770 1.260 0.790 2.660 ;
        RECT  0.790 1.260 1.190 3.150 ;
        RECT  1.190 1.260 1.210 2.660 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.180 5.440 ;
        RECT  0.180 4.010 0.580 5.440 ;
        RECT  0.580 4.640 1.420 5.440 ;
        RECT  1.420 4.010 1.820 5.440 ;
        RECT  1.820 4.640 3.500 5.440 ;
        RECT  3.500 4.070 3.900 5.440 ;
        RECT  3.900 4.640 5.960 5.440 ;
        RECT  5.960 3.990 6.360 5.440 ;
        RECT  6.360 4.640 8.420 5.440 ;
        RECT  8.420 3.970 8.820 5.440 ;
        RECT  8.820 4.640 10.300 5.440 ;
        RECT  10.300 3.960 10.700 5.440 ;
        RECT  10.700 4.640 11.970 5.440 ;
        RECT  11.970 3.960 12.370 5.440 ;
        RECT  12.370 4.640 12.540 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.990 ;
        RECT  0.570 -0.400 1.410 0.400 ;
        RECT  1.410 -0.400 1.810 0.990 ;
        RECT  1.810 -0.400 3.030 0.400 ;
        RECT  3.030 -0.400 3.430 0.560 ;
        RECT  3.430 -0.400 4.490 0.400 ;
        RECT  4.490 -0.400 4.890 0.560 ;
        RECT  4.890 -0.400 5.950 0.400 ;
        RECT  5.950 -0.400 6.350 0.560 ;
        RECT  6.350 -0.400 7.410 0.400 ;
        RECT  7.410 -0.400 7.810 0.560 ;
        RECT  7.810 -0.400 8.870 0.400 ;
        RECT  8.870 -0.400 9.270 0.560 ;
        RECT  9.270 -0.400 10.460 0.400 ;
        RECT  10.460 -0.400 10.860 0.990 ;
        RECT  10.860 -0.400 11.880 0.400 ;
        RECT  11.880 -0.400 12.280 0.990 ;
        RECT  12.280 -0.400 12.540 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.040 2.180 12.280 3.670 ;
        RECT  9.080 3.430 12.040 3.670 ;
        RECT  9.720 1.030 10.010 1.430 ;
        RECT  9.720 2.750 9.880 3.150 ;
        RECT  9.480 1.030 9.720 3.150 ;
        RECT  9.360 1.850 9.480 2.250 ;
        RECT  8.840 1.300 9.080 3.670 ;
        RECT  8.540 1.300 8.840 1.540 ;
        RECT  7.600 3.210 8.840 3.670 ;
        RECT  8.170 2.260 8.570 2.660 ;
        RECT  8.140 1.220 8.540 1.620 ;
        RECT  6.470 2.340 8.170 2.580 ;
        RECT  7.080 1.300 8.140 1.540 ;
        RECT  7.200 3.210 7.600 4.190 ;
        RECT  6.920 1.220 7.080 1.620 ;
        RECT  6.680 1.220 6.920 2.060 ;
        RECT  5.850 1.820 6.680 2.060 ;
        RECT  6.230 2.340 6.470 3.450 ;
        RECT  5.120 3.210 6.230 3.450 ;
        RECT  5.610 1.820 5.850 2.500 ;
        RECT  4.160 1.300 5.620 1.540 ;
        RECT  4.070 2.260 5.610 2.500 ;
        RECT  4.720 3.210 5.120 4.190 ;
        RECT  3.560 3.210 4.720 3.670 ;
        RECT  3.760 1.220 4.160 1.620 ;
        RECT  3.830 2.260 4.070 2.660 ;
        RECT  3.560 1.380 3.760 1.620 ;
        RECT  3.320 1.380 3.560 3.670 ;
        RECT  0.500 3.430 3.320 3.670 ;
        RECT  2.800 1.310 3.040 2.990 ;
        RECT  2.610 1.310 2.800 1.550 ;
        RECT  2.710 2.750 2.800 2.990 ;
        RECT  2.310 2.750 2.710 3.150 ;
        RECT  2.210 1.150 2.610 1.550 ;
        RECT  0.260 2.180 0.500 3.670 ;
    END
END RSLATNX4

MACRO RSLATNX2
    CLASS CORE ;
    FOREIGN RSLATNX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ RSLATNXL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.410 2.160 3.760 2.760 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 1.830 4.230 2.090 ;
        RECT  4.230 1.690 4.630 2.090 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.800 2.950 6.910 3.210 ;
        RECT  6.910 2.950 7.350 3.220 ;
        RECT  7.350 2.950 7.510 3.990 ;
        RECT  7.350 1.000 7.510 1.400 ;
        RECT  7.510 1.000 7.750 3.990 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.160 0.890 0.170 4.100 ;
        RECT  0.170 0.890 0.400 4.110 ;
        RECT  0.400 3.130 0.570 4.110 ;
        RECT  0.400 0.890 0.570 1.290 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.920 5.440 ;
        RECT  0.920 4.090 0.930 5.440 ;
        RECT  0.930 3.890 1.330 5.440 ;
        RECT  1.330 4.090 1.340 5.440 ;
        RECT  1.340 4.640 3.740 5.440 ;
        RECT  3.740 4.480 4.140 5.440 ;
        RECT  4.140 4.640 6.500 5.440 ;
        RECT  6.500 4.370 6.510 5.440 ;
        RECT  6.510 4.170 6.910 5.440 ;
        RECT  6.910 4.370 6.920 5.440 ;
        RECT  6.920 4.640 7.920 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.920 0.400 ;
        RECT  0.920 -0.400 0.930 1.130 ;
        RECT  0.930 -0.400 1.330 1.330 ;
        RECT  1.330 -0.400 1.340 1.130 ;
        RECT  1.340 -0.400 2.440 0.400 ;
        RECT  2.440 -0.400 2.450 1.130 ;
        RECT  2.450 -0.400 2.850 1.330 ;
        RECT  2.850 -0.400 2.860 1.130 ;
        RECT  2.860 -0.400 5.010 0.400 ;
        RECT  5.010 -0.400 5.410 0.560 ;
        RECT  5.410 -0.400 6.580 0.400 ;
        RECT  6.580 -0.400 6.590 1.130 ;
        RECT  6.590 -0.400 6.990 1.330 ;
        RECT  6.990 -0.400 7.000 1.130 ;
        RECT  7.000 -0.400 7.920 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.990 1.720 7.230 2.370 ;
        RECT  6.230 1.720 6.990 1.960 ;
        RECT  6.430 2.260 6.590 2.660 ;
        RECT  6.190 2.260 6.430 3.890 ;
        RECT  5.910 1.300 6.230 1.960 ;
        RECT  6.130 3.650 6.190 3.890 ;
        RECT  5.890 3.650 6.130 4.180 ;
        RECT  5.830 1.300 5.910 3.350 ;
        RECT  2.100 3.940 5.890 4.180 ;
        RECT  5.670 1.720 5.830 3.350 ;
        RECT  5.610 3.110 5.670 3.350 ;
        RECT  5.370 3.110 5.610 3.660 ;
        RECT  5.150 1.170 5.390 2.660 ;
        RECT  2.620 3.420 5.370 3.660 ;
        RECT  4.130 1.170 5.150 1.410 ;
        RECT  4.870 2.420 5.150 2.660 ;
        RECT  4.630 2.420 4.870 3.140 ;
        RECT  4.470 2.740 4.630 3.140 ;
        RECT  3.330 1.370 3.730 1.850 ;
        RECT  3.140 1.610 3.330 1.850 ;
        RECT  2.900 1.610 3.140 3.140 ;
        RECT  2.040 2.170 2.900 2.570 ;
        RECT  2.380 2.850 2.620 3.660 ;
        RECT  1.640 2.850 2.380 3.090 ;
        RECT  1.860 3.370 2.100 4.180 ;
        RECT  1.690 1.260 2.090 1.870 ;
        RECT  1.120 3.370 1.860 3.610 ;
        RECT  1.120 1.630 1.690 1.870 ;
        RECT  1.400 2.170 1.640 3.090 ;
        RECT  0.880 1.630 1.120 3.610 ;
        RECT  0.680 2.170 0.880 2.590 ;
    END
END RSLATNX2

MACRO RSLATNX1
    CLASS CORE ;
    FOREIGN RSLATNX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ RSLATNXL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.070 2.370 3.410 2.610 ;
        RECT  3.410 1.850 3.500 2.610 ;
        RECT  3.500 1.830 3.650 2.610 ;
        RECT  3.650 1.830 3.760 2.090 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.910 2.370 4.510 2.670 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.140 2.950 6.150 3.210 ;
        RECT  6.150 2.870 6.810 3.270 ;
        RECT  6.690 1.390 6.810 1.790 ;
        RECT  6.810 2.640 6.850 3.270 ;
        RECT  6.810 1.390 6.850 1.840 ;
        RECT  6.850 1.390 7.090 3.270 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.160 3.510 0.170 4.130 ;
        RECT  0.170 1.390 0.410 4.130 ;
        RECT  0.410 1.390 0.450 1.840 ;
        RECT  0.450 1.390 0.570 1.790 ;
        RECT  0.410 3.510 0.580 4.130 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.980 5.440 ;
        RECT  0.980 3.900 0.990 5.440 ;
        RECT  0.990 3.700 1.390 5.440 ;
        RECT  1.390 3.900 1.400 5.440 ;
        RECT  1.400 4.640 3.250 5.440 ;
        RECT  3.250 4.480 3.650 5.440 ;
        RECT  3.650 4.640 6.080 5.440 ;
        RECT  6.080 4.480 6.480 5.440 ;
        RECT  6.480 4.640 7.260 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.910 0.400 ;
        RECT  0.910 -0.400 1.310 0.560 ;
        RECT  1.310 -0.400 2.720 0.400 ;
        RECT  2.720 -0.400 3.120 0.560 ;
        RECT  3.120 -0.400 4.390 0.400 ;
        RECT  4.390 -0.400 4.790 0.560 ;
        RECT  4.790 -0.400 6.530 0.400 ;
        RECT  6.530 -0.400 6.930 0.560 ;
        RECT  6.930 -0.400 7.260 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.250 2.090 6.570 2.490 ;
        RECT  6.010 0.800 6.250 2.490 ;
        RECT  5.610 0.800 6.010 1.040 ;
        RECT  5.760 2.250 6.010 2.490 ;
        RECT  5.520 2.250 5.760 3.850 ;
        RECT  5.490 1.330 5.730 1.810 ;
        RECT  5.370 0.720 5.610 1.040 ;
        RECT  5.210 3.610 5.520 3.850 ;
        RECT  4.930 1.330 5.490 1.570 ;
        RECT  5.210 0.720 5.370 0.960 ;
        RECT  5.020 2.430 5.210 2.830 ;
        RECT  4.810 3.610 5.210 4.010 ;
        RECT  4.780 1.850 5.020 3.190 ;
        RECT  4.690 0.860 4.930 1.570 ;
        RECT  2.870 3.770 4.810 4.010 ;
        RECT  4.410 1.850 4.780 2.090 ;
        RECT  4.290 2.950 4.780 3.190 ;
        RECT  2.130 0.860 4.690 1.100 ;
        RECT  4.170 1.380 4.410 2.090 ;
        RECT  2.790 2.940 3.850 3.180 ;
        RECT  2.790 1.380 2.870 1.790 ;
        RECT  2.630 3.770 2.870 4.370 ;
        RECT  2.630 1.380 2.790 3.180 ;
        RECT  2.550 1.550 2.630 3.180 ;
        RECT  2.470 4.130 2.630 4.370 ;
        RECT  1.370 1.550 2.550 1.950 ;
        RECT  1.730 0.720 2.130 1.100 ;
        RECT  1.510 2.910 1.910 3.310 ;
        RECT  1.090 0.860 1.730 1.100 ;
        RECT  1.090 2.910 1.510 3.150 ;
        RECT  0.850 0.860 1.090 3.150 ;
        RECT  0.730 2.070 0.850 2.470 ;
    END
END RSLATNX1

MACRO RSLATXL
    CLASS CORE ;
    FOREIGN RSLATXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 1.820 3.200 2.360 ;
        END
    END S
    PIN R
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.860 2.380 4.510 2.720 ;
        END
    END R
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.170 1.190 0.410 3.540 ;
        RECT  0.410 2.950 0.570 3.540 ;
        RECT  0.410 1.190 0.570 1.590 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.140 3.510 6.150 3.770 ;
        RECT  6.690 1.280 6.810 1.680 ;
        RECT  6.150 3.510 6.850 3.910 ;
        RECT  6.810 1.280 6.850 1.840 ;
        RECT  6.850 1.280 7.090 3.910 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.950 5.440 ;
        RECT  0.950 4.480 1.030 5.440 ;
        RECT  1.030 4.460 2.110 5.440 ;
        RECT  2.110 4.480 2.480 5.440 ;
        RECT  2.480 4.640 4.960 5.440 ;
        RECT  4.960 4.480 5.940 5.440 ;
        RECT  5.940 4.640 7.260 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.850 0.400 ;
        RECT  0.850 -0.400 1.250 0.560 ;
        RECT  1.250 -0.400 2.970 0.400 ;
        RECT  2.970 -0.400 3.370 0.560 ;
        RECT  3.370 -0.400 6.030 0.400 ;
        RECT  6.030 -0.400 6.430 0.560 ;
        RECT  6.430 -0.400 7.260 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.700 2.090 6.550 2.490 ;
        RECT  5.460 1.350 5.700 3.750 ;
        RECT  4.690 1.350 5.460 1.590 ;
        RECT  4.690 3.510 5.460 3.750 ;
        RECT  5.020 2.580 5.180 2.980 ;
        RECT  4.780 1.870 5.020 3.230 ;
        RECT  3.890 0.730 4.950 0.970 ;
        RECT  4.330 1.870 4.780 2.110 ;
        RECT  4.170 2.990 4.780 3.230 ;
        RECT  4.450 3.510 4.690 4.360 ;
        RECT  2.990 4.120 4.450 4.360 ;
        RECT  4.090 1.460 4.330 2.110 ;
        RECT  3.930 2.990 4.170 3.840 ;
        RECT  3.930 1.460 4.090 1.700 ;
        RECT  3.270 3.600 3.930 3.840 ;
        RECT  3.650 0.730 3.890 1.100 ;
        RECT  2.690 0.860 3.650 1.100 ;
        RECT  2.570 2.860 3.590 3.100 ;
        RECT  2.750 3.660 2.990 4.360 ;
        RECT  1.350 3.660 2.750 3.900 ;
        RECT  2.450 0.670 2.690 1.100 ;
        RECT  2.480 2.370 2.570 3.100 ;
        RECT  2.330 1.380 2.480 3.100 ;
        RECT  1.830 0.670 2.450 0.910 ;
        RECT  2.240 1.380 2.330 2.620 ;
        RECT  1.950 2.220 2.240 2.620 ;
        RECT  1.270 2.980 2.050 3.220 ;
        RECT  1.590 0.670 1.830 1.210 ;
        RECT  1.270 0.970 1.590 1.210 ;
        RECT  1.030 0.970 1.270 3.220 ;
        RECT  0.690 1.870 1.030 2.110 ;
    END
END RSLATXL

MACRO RSLATX4
    CLASS CORE ;
    FOREIGN RSLATX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ RSLATXL ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.940 1.760 10.500 2.170 ;
        END
    END S
    PIN R
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 1.830 2.440 2.090 ;
        RECT  2.440 1.850 2.460 2.090 ;
        RECT  2.460 1.850 2.860 2.350 ;
        END
    END R
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.330 1.820 11.350 3.220 ;
        RECT  11.350 1.430 11.360 3.220 ;
        RECT  11.360 1.230 11.760 3.220 ;
        RECT  11.760 1.430 11.770 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.770 1.820 0.780 3.220 ;
        RECT  0.780 1.370 0.870 3.220 ;
        RECT  0.870 1.370 1.190 3.450 ;
        RECT  1.190 1.370 1.210 3.610 ;
        RECT  1.210 1.370 1.470 1.790 ;
        RECT  1.210 3.210 1.590 3.610 ;
        RECT  1.470 1.380 1.670 1.780 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.560 5.440 ;
        RECT  0.560 4.210 0.570 5.440 ;
        RECT  0.570 4.010 0.970 5.440 ;
        RECT  0.970 4.210 0.980 5.440 ;
        RECT  0.980 4.640 1.870 5.440 ;
        RECT  1.870 4.210 1.880 5.440 ;
        RECT  1.880 4.010 2.280 5.440 ;
        RECT  2.280 4.210 2.290 5.440 ;
        RECT  2.290 4.640 3.440 5.440 ;
        RECT  3.440 4.480 3.840 5.440 ;
        RECT  3.840 4.640 5.030 5.440 ;
        RECT  5.030 3.730 5.040 5.440 ;
        RECT  5.040 3.530 5.440 5.440 ;
        RECT  5.440 3.730 5.450 5.440 ;
        RECT  5.450 4.640 6.330 5.440 ;
        RECT  6.330 3.730 6.340 5.440 ;
        RECT  6.340 3.530 6.740 5.440 ;
        RECT  6.740 3.730 6.750 5.440 ;
        RECT  6.750 4.640 7.730 5.440 ;
        RECT  7.730 3.730 7.740 5.440 ;
        RECT  7.740 3.530 8.140 5.440 ;
        RECT  8.140 3.730 8.150 5.440 ;
        RECT  8.150 4.640 9.080 5.440 ;
        RECT  9.080 4.480 9.480 5.440 ;
        RECT  9.480 4.640 10.710 5.440 ;
        RECT  10.710 4.250 10.720 5.440 ;
        RECT  10.720 4.130 11.120 5.440 ;
        RECT  11.120 4.250 11.130 5.440 ;
        RECT  11.130 4.640 11.960 5.440 ;
        RECT  11.960 4.250 11.970 5.440 ;
        RECT  11.970 4.130 12.370 5.440 ;
        RECT  12.370 4.250 12.380 5.440 ;
        RECT  12.380 4.640 12.540 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.590 0.400 ;
        RECT  0.590 -0.400 0.600 0.900 ;
        RECT  0.600 -0.400 1.000 1.100 ;
        RECT  1.000 -0.400 1.010 0.900 ;
        RECT  1.010 -0.400 1.870 0.400 ;
        RECT  1.870 -0.400 1.880 0.900 ;
        RECT  1.880 -0.400 2.280 1.100 ;
        RECT  2.280 -0.400 2.290 0.900 ;
        RECT  2.290 -0.400 3.980 0.400 ;
        RECT  3.980 -0.400 3.990 0.670 ;
        RECT  3.990 -0.400 4.390 0.870 ;
        RECT  4.390 -0.400 4.400 0.670 ;
        RECT  4.400 -0.400 6.420 0.400 ;
        RECT  6.420 -0.400 6.430 0.670 ;
        RECT  6.430 -0.400 6.830 0.870 ;
        RECT  6.830 -0.400 6.840 0.670 ;
        RECT  6.840 -0.400 9.070 0.400 ;
        RECT  9.070 -0.400 9.470 0.560 ;
        RECT  9.470 -0.400 10.680 0.400 ;
        RECT  10.680 -0.400 10.690 0.750 ;
        RECT  10.690 -0.400 11.090 0.950 ;
        RECT  11.090 -0.400 11.100 0.750 ;
        RECT  11.100 -0.400 11.960 0.400 ;
        RECT  11.960 -0.400 11.970 0.750 ;
        RECT  11.970 -0.400 12.370 0.950 ;
        RECT  12.370 -0.400 12.380 0.750 ;
        RECT  12.380 -0.400 12.540 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.040 2.120 12.280 3.850 ;
        RECT  8.920 3.610 12.040 3.850 ;
        RECT  10.760 1.230 11.000 3.330 ;
        RECT  10.260 1.230 10.760 1.470 ;
        RECT  9.910 3.090 10.760 3.330 ;
        RECT  10.020 0.690 10.260 1.470 ;
        RECT  9.860 0.690 10.020 1.090 ;
        RECT  9.670 2.440 9.910 3.330 ;
        RECT  9.510 2.440 9.670 2.840 ;
        RECT  8.760 1.720 9.160 2.120 ;
        RECT  8.680 2.750 8.920 3.850 ;
        RECT  8.750 1.720 8.760 1.960 ;
        RECT  8.510 0.670 8.750 1.960 ;
        RECT  8.410 2.750 8.680 3.150 ;
        RECT  7.450 0.670 8.510 0.910 ;
        RECT  8.130 2.750 8.410 3.020 ;
        RECT  7.730 1.190 8.130 3.020 ;
        RECT  7.410 2.780 7.730 3.020 ;
        RECT  7.210 0.670 7.450 2.470 ;
        RECT  7.010 2.780 7.410 3.180 ;
        RECT  7.050 1.150 7.210 2.470 ;
        RECT  5.610 1.150 7.050 1.390 ;
        RECT  6.710 2.780 7.010 3.020 ;
        RECT  6.470 2.310 6.710 3.020 ;
        RECT  6.380 2.310 6.470 2.550 ;
        RECT  5.980 2.150 6.380 2.550 ;
        RECT  5.700 2.850 6.100 3.250 ;
        RECT  4.570 2.310 5.980 2.550 ;
        RECT  4.610 3.010 5.700 3.250 ;
        RECT  5.210 0.940 5.610 1.390 ;
        RECT  4.050 1.150 5.210 1.390 ;
        RECT  4.050 3.010 4.610 3.410 ;
        RECT  4.330 1.720 4.570 2.550 ;
        RECT  3.810 1.150 4.050 3.730 ;
        RECT  2.200 3.490 3.810 3.730 ;
        RECT  3.290 1.150 3.530 3.210 ;
        RECT  2.700 1.150 3.290 1.390 ;
        RECT  2.680 2.970 3.290 3.210 ;
        RECT  1.960 2.680 2.200 3.730 ;
        RECT  1.820 2.680 1.960 2.920 ;
        RECT  1.580 2.180 1.820 2.920 ;
    END
END RSLATX4

MACRO RSLATX2
    CLASS CORE ;
    FOREIGN RSLATX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ RSLATXL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.140 2.390 6.150 2.650 ;
        RECT  6.150 2.070 6.400 2.650 ;
        RECT  6.400 2.070 6.590 2.470 ;
        END
    END S
    PIN R
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 0.870 3.210 ;
        RECT  0.870 2.750 1.120 3.210 ;
        RECT  1.120 2.750 1.260 2.990 ;
        RECT  1.260 2.590 1.660 2.990 ;
        END
    END R
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  7.350 3.130 7.520 4.110 ;
        RECT  7.430 0.700 7.520 1.680 ;
        RECT  7.520 0.700 7.670 4.110 ;
        RECT  7.670 0.710 7.750 4.110 ;
        RECT  7.750 0.710 7.760 4.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.210 2.090 ;
        RECT  0.210 0.670 0.250 4.090 ;
        RECT  0.250 0.660 0.450 4.100 ;
        RECT  0.450 0.660 0.460 2.090 ;
        RECT  0.450 3.120 0.490 4.100 ;
        RECT  0.460 0.660 0.490 1.860 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 4.480 2.160 5.440 ;
        RECT  2.160 4.640 3.880 5.440 ;
        RECT  3.880 4.480 4.280 5.440 ;
        RECT  4.280 4.640 5.450 5.440 ;
        RECT  5.450 3.790 5.460 5.440 ;
        RECT  5.460 3.590 5.860 5.440 ;
        RECT  5.860 3.790 5.870 5.440 ;
        RECT  5.870 4.640 6.580 5.440 ;
        RECT  6.580 3.980 6.590 5.440 ;
        RECT  6.590 3.780 6.990 5.440 ;
        RECT  6.990 3.980 7.000 5.440 ;
        RECT  7.000 4.640 7.920 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        RECT  0.990 -0.400 1.390 0.560 ;
        RECT  1.390 -0.400 2.200 0.400 ;
        RECT  2.200 -0.400 2.600 0.560 ;
        RECT  2.600 -0.400 4.110 0.400 ;
        RECT  4.110 -0.400 4.510 0.560 ;
        RECT  4.510 -0.400 6.530 0.400 ;
        RECT  6.530 -0.400 6.930 0.560 ;
        RECT  6.930 -0.400 7.920 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  7.150 1.950 7.280 2.350 ;
        RECT  6.910 0.860 7.150 2.350 ;
        RECT  5.790 0.860 6.910 1.100 ;
        RECT  5.710 2.930 6.360 3.170 ;
        RECT  5.710 1.460 6.290 1.700 ;
        RECT  5.390 0.720 5.790 1.100 ;
        RECT  5.470 1.460 5.710 3.170 ;
        RECT  5.180 0.860 5.390 1.100 ;
        RECT  4.940 0.860 5.180 3.880 ;
        RECT  4.700 3.480 4.940 3.880 ;
        RECT  2.780 3.640 4.700 3.880 ;
        RECT  4.500 2.020 4.660 2.420 ;
        RECT  4.260 1.080 4.500 3.190 ;
        RECT  2.720 1.080 4.260 1.320 ;
        RECT  3.550 2.950 4.260 3.190 ;
        RECT  3.350 1.650 3.750 2.200 ;
        RECT  3.150 2.950 3.550 3.350 ;
        RECT  2.180 1.650 3.350 1.890 ;
        RECT  2.780 2.170 2.860 2.570 ;
        RECT  2.540 2.170 2.780 3.880 ;
        RECT  2.480 0.860 2.720 1.320 ;
        RECT  2.460 2.170 2.540 2.570 ;
        RECT  1.060 0.860 2.480 1.100 ;
        RECT  1.940 1.380 2.180 3.670 ;
        RECT  1.760 1.380 1.940 1.780 ;
        RECT  1.700 3.270 1.940 3.670 ;
        RECT  0.820 0.860 1.060 2.270 ;
    END
END RSLATX2

MACRO RSLATX1
    CLASS CORE ;
    FOREIGN RSLATX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ RSLATXL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.750 1.820 3.100 2.480 ;
        END
    END S
    PIN R
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.660 2.380 4.510 2.720 ;
        END
    END R
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.160 1.080 0.400 3.770 ;
        RECT  0.400 3.040 0.460 3.770 ;
        RECT  0.460 3.040 0.550 3.500 ;
        RECT  0.550 3.040 0.570 3.440 ;
        RECT  0.400 1.080 0.570 1.480 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.140 2.950 6.580 3.220 ;
        RECT  6.580 1.320 6.710 1.720 ;
        RECT  6.580 2.950 6.740 3.670 ;
        RECT  6.710 1.320 6.740 1.820 ;
        RECT  6.740 1.320 6.980 3.670 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.370 5.440 ;
        RECT  1.370 4.480 1.450 5.440 ;
        RECT  1.450 4.460 2.250 5.440 ;
        RECT  2.250 4.480 2.330 5.440 ;
        RECT  2.330 4.640 4.790 5.440 ;
        RECT  4.790 4.480 4.870 5.440 ;
        RECT  4.870 4.460 5.670 5.440 ;
        RECT  5.670 4.480 5.750 5.440 ;
        RECT  5.750 4.640 7.260 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.790 0.400 ;
        RECT  0.790 -0.400 1.190 0.560 ;
        RECT  1.190 -0.400 2.850 0.400 ;
        RECT  2.850 -0.400 3.250 0.560 ;
        RECT  3.250 -0.400 5.750 0.400 ;
        RECT  5.750 -0.400 6.150 0.560 ;
        RECT  6.150 -0.400 7.260 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.780 2.090 6.460 2.490 ;
        RECT  5.540 1.350 5.780 3.810 ;
        RECT  4.470 1.350 5.540 1.590 ;
        RECT  4.510 3.570 5.540 3.810 ;
        RECT  4.790 1.870 5.030 3.290 ;
        RECT  4.130 1.870 4.790 2.110 ;
        RECT  3.990 3.050 4.790 3.290 ;
        RECT  4.190 0.730 4.670 0.970 ;
        RECT  4.270 3.570 4.510 4.360 ;
        RECT  2.850 4.120 4.270 4.360 ;
        RECT  3.950 0.730 4.190 1.100 ;
        RECT  3.890 1.380 4.130 2.110 ;
        RECT  3.750 3.050 3.990 3.840 ;
        RECT  2.490 0.860 3.950 1.100 ;
        RECT  3.730 1.380 3.890 1.780 ;
        RECT  3.150 3.600 3.750 3.840 ;
        RECT  3.150 2.750 3.390 3.180 ;
        RECT  2.450 2.750 3.150 2.990 ;
        RECT  2.610 3.660 2.850 4.360 ;
        RECT  1.350 3.660 2.610 3.900 ;
        RECT  2.090 0.670 2.490 1.100 ;
        RECT  2.210 1.380 2.450 2.990 ;
        RECT  1.980 2.080 2.210 2.480 ;
        RECT  1.690 0.860 2.090 1.100 ;
        RECT  1.690 2.760 1.910 3.290 ;
        RECT  1.670 0.860 1.690 3.290 ;
        RECT  1.450 0.860 1.670 3.000 ;
        RECT  0.900 1.760 1.450 2.180 ;
        RECT  0.750 1.770 0.900 2.170 ;
    END
END RSLATX1

MACRO OR4XL
    CLASS CORE ;
    FOREIGN OR4XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.630 2.950 4.170 3.350 ;
        RECT  4.160 1.830 4.170 2.090 ;
        RECT  4.050 0.900 4.170 1.300 ;
        RECT  4.170 0.900 4.290 3.350 ;
        RECT  4.290 0.900 4.410 3.190 ;
        RECT  4.410 1.830 4.420 2.090 ;
        RECT  4.410 0.900 4.450 1.300 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.530 2.360 3.100 2.800 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.010 1.590 2.020 1.830 ;
        RECT  2.020 1.590 2.430 2.090 ;
        RECT  2.430 1.830 2.440 2.090 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.350 1.740 1.590 2.650 ;
        RECT  1.590 2.390 1.780 2.650 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.060 0.550 2.690 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 2.750 5.440 ;
        RECT  2.750 4.480 3.150 5.440 ;
        RECT  3.150 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.500 0.400 ;
        RECT  1.500 -0.400 1.900 0.560 ;
        RECT  1.900 -0.400 3.180 0.400 ;
        RECT  3.180 -0.400 3.580 0.560 ;
        RECT  3.580 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.630 1.580 3.800 1.980 ;
        RECT  3.400 1.070 3.630 1.980 ;
        RECT  3.390 1.070 3.400 1.900 ;
        RECT  2.770 1.070 3.390 1.310 ;
        RECT  2.370 0.910 2.770 1.310 ;
        RECT  1.230 1.070 2.370 1.310 ;
        RECT  1.070 1.050 1.230 1.450 ;
        RECT  0.830 1.050 1.070 3.360 ;
        RECT  0.550 2.960 0.830 3.360 ;
    END
END OR4XL

MACRO OR4X4
    CLASS CORE ;
    FOREIGN OR4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OR4XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  5.390 1.820 5.410 3.220 ;
        RECT  5.410 1.350 5.830 3.220 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.430 2.310 0.770 2.710 ;
        RECT  0.770 2.310 0.780 3.100 ;
        RECT  0.780 2.310 0.860 3.760 ;
        RECT  0.860 2.310 1.020 3.770 ;
        RECT  1.020 3.510 1.120 3.770 ;
        RECT  1.120 3.520 3.460 3.760 ;
        RECT  3.460 2.920 3.700 3.760 ;
        RECT  3.700 2.920 4.330 3.160 ;
        RECT  4.330 2.760 4.570 3.160 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.560 1.410 0.960 1.990 ;
        RECT  0.960 1.410 3.770 1.650 ;
        RECT  3.770 1.410 4.010 2.440 ;
        RECT  4.010 1.820 4.200 2.440 ;
        RECT  4.200 1.820 4.310 2.090 ;
        RECT  4.310 1.830 4.420 2.090 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.390 1.600 2.650 ;
        RECT  1.600 1.930 1.780 2.650 ;
        RECT  1.780 1.930 1.870 2.630 ;
        RECT  1.870 1.930 2.000 2.330 ;
        RECT  2.000 1.930 3.090 2.170 ;
        RECT  3.090 1.930 3.490 2.440 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.370 2.450 2.770 3.190 ;
        RECT  2.770 2.950 2.840 3.190 ;
        RECT  2.840 2.950 3.100 3.210 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.250 5.440 ;
        RECT  0.250 3.180 0.490 5.440 ;
        RECT  0.490 4.640 4.620 5.440 ;
        RECT  4.620 4.210 4.630 5.440 ;
        RECT  4.630 4.010 5.030 5.440 ;
        RECT  5.030 4.210 5.040 5.440 ;
        RECT  5.040 4.640 6.020 5.440 ;
        RECT  6.020 4.210 6.030 5.440 ;
        RECT  6.030 4.010 6.430 5.440 ;
        RECT  6.430 4.210 6.440 5.440 ;
        RECT  6.440 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.050 0.400 ;
        RECT  1.050 -0.400 1.450 0.560 ;
        RECT  1.450 -0.400 3.250 0.400 ;
        RECT  3.250 -0.400 3.650 0.560 ;
        RECT  3.650 -0.400 4.780 0.400 ;
        RECT  4.780 -0.400 4.790 0.870 ;
        RECT  4.790 -0.400 5.190 0.990 ;
        RECT  5.190 -0.400 5.200 0.870 ;
        RECT  5.200 -0.400 6.020 0.400 ;
        RECT  6.020 -0.400 6.030 0.870 ;
        RECT  6.030 -0.400 6.430 1.070 ;
        RECT  6.430 -0.400 6.440 0.870 ;
        RECT  6.440 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.100 2.180 6.340 3.730 ;
        RECT  5.090 3.490 6.100 3.730 ;
        RECT  4.850 1.310 5.090 3.730 ;
        RECT  4.530 1.310 4.850 1.550 ;
        RECT  4.220 3.490 4.850 3.730 ;
        RECT  4.290 0.890 4.530 1.550 ;
        RECT  0.230 0.890 4.290 1.130 ;
        RECT  3.980 3.490 4.220 4.280 ;
        RECT  2.370 4.040 3.980 4.280 ;
    END
END OR4X4

MACRO OR4X2
    CLASS CORE ;
    FOREIGN OR4X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OR4XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.040 0.790 4.050 1.350 ;
        RECT  3.820 3.210 4.170 4.190 ;
        RECT  4.160 1.830 4.170 2.090 ;
        RECT  4.050 0.670 4.170 1.550 ;
        RECT  4.170 0.670 4.220 4.190 ;
        RECT  4.220 0.670 4.410 4.180 ;
        RECT  4.410 1.830 4.420 2.090 ;
        RECT  4.410 0.670 4.450 1.550 ;
        RECT  4.450 0.790 4.460 1.350 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.530 2.360 3.100 2.780 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.000 1.620 2.440 2.100 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.370 1.860 1.610 2.650 ;
        RECT  1.610 2.390 1.780 2.650 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.060 0.550 2.710 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 2.840 5.440 ;
        RECT  2.840 4.480 3.240 5.440 ;
        RECT  3.240 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.620 0.400 ;
        RECT  1.620 -0.400 2.020 0.560 ;
        RECT  2.020 -0.400 3.220 0.400 ;
        RECT  3.220 -0.400 3.230 0.410 ;
        RECT  3.230 -0.400 3.630 0.560 ;
        RECT  3.630 -0.400 3.640 0.410 ;
        RECT  3.640 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.630 1.780 3.800 2.180 ;
        RECT  3.400 1.110 3.630 2.180 ;
        RECT  3.390 1.110 3.400 2.100 ;
        RECT  2.770 1.110 3.390 1.350 ;
        RECT  2.370 0.950 2.770 1.350 ;
        RECT  1.230 1.110 2.370 1.350 ;
        RECT  1.060 1.050 1.230 1.450 ;
        RECT  0.830 1.050 1.060 3.680 ;
        RECT  0.820 1.060 0.830 3.680 ;
        RECT  0.550 3.280 0.820 3.680 ;
    END
END OR4X2

MACRO OR4X1
    CLASS CORE ;
    FOREIGN OR4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OR4XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.630 3.080 4.170 3.480 ;
        RECT  4.160 1.830 4.170 2.090 ;
        RECT  4.050 1.030 4.170 1.430 ;
        RECT  4.170 1.030 4.410 3.480 ;
        RECT  4.410 1.830 4.420 2.090 ;
        RECT  4.410 1.030 4.450 1.430 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.530 2.360 3.100 2.800 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.000 1.760 2.010 2.090 ;
        RECT  2.010 1.590 2.430 2.090 ;
        RECT  2.430 1.830 2.440 2.090 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.370 1.860 1.610 2.650 ;
        RECT  1.610 2.390 1.780 2.650 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.060 0.460 2.650 ;
        RECT  0.460 2.060 0.540 2.640 ;
        RECT  0.540 2.060 0.550 2.440 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 2.770 5.440 ;
        RECT  2.770 4.480 3.170 5.440 ;
        RECT  3.170 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.620 0.400 ;
        RECT  1.620 -0.400 2.020 0.560 ;
        RECT  2.020 -0.400 3.240 0.400 ;
        RECT  3.240 -0.400 3.640 0.560 ;
        RECT  3.640 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.620 1.700 3.790 2.100 ;
        RECT  3.390 1.070 3.620 2.100 ;
        RECT  3.380 1.070 3.390 2.020 ;
        RECT  2.770 1.070 3.380 1.310 ;
        RECT  2.370 0.910 2.770 1.310 ;
        RECT  1.230 1.050 2.370 1.290 ;
        RECT  1.060 1.050 1.230 1.450 ;
        RECT  0.830 1.050 1.060 3.360 ;
        RECT  0.820 1.060 0.830 3.360 ;
        RECT  0.570 2.960 0.820 3.360 ;
    END
END OR4X1

MACRO OR3XL
    CLASS CORE ;
    FOREIGN OR3XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.160 2.950 3.510 3.350 ;
        RECT  3.500 1.830 3.510 2.090 ;
        RECT  3.390 1.020 3.510 1.420 ;
        RECT  3.510 1.020 3.750 3.350 ;
        RECT  3.750 1.830 3.760 2.090 ;
        RECT  3.750 1.020 3.790 1.420 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.870 2.360 2.440 2.800 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.400 1.580 1.870 2.100 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.310 0.690 2.650 ;
        RECT  0.690 2.230 1.090 2.650 ;
        RECT  1.090 2.390 1.120 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 2.180 5.440 ;
        RECT  2.180 4.480 2.580 5.440 ;
        RECT  2.580 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.960 0.400 ;
        RECT  0.960 -0.400 1.360 0.560 ;
        RECT  1.360 -0.400 2.560 0.400 ;
        RECT  2.560 -0.400 2.570 0.410 ;
        RECT  2.570 -0.400 2.970 0.560 ;
        RECT  2.970 -0.400 2.980 0.410 ;
        RECT  2.980 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.980 1.700 3.140 2.100 ;
        RECT  2.740 1.070 2.980 2.100 ;
        RECT  2.110 1.070 2.740 1.310 ;
        RECT  1.710 0.910 2.110 1.310 ;
        RECT  0.580 1.070 1.710 1.310 ;
        RECT  0.420 2.960 0.750 3.360 ;
        RECT  0.420 0.910 0.580 1.310 ;
        RECT  0.180 0.910 0.420 3.360 ;
    END
END OR3XL

MACRO OR3X4
    CLASS CORE ;
    FOREIGN OR3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OR3XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.730 1.260 4.750 2.660 ;
        RECT  4.750 1.260 4.760 3.080 ;
        RECT  4.760 1.150 5.160 3.150 ;
        RECT  5.160 1.260 5.170 3.090 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.690 1.790 0.770 2.210 ;
        RECT  0.770 1.790 1.120 2.220 ;
        RECT  1.120 1.790 3.380 2.030 ;
        RECT  3.380 1.670 3.780 2.030 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 2.310 1.520 2.640 ;
        RECT  1.520 2.310 1.780 2.650 ;
        RECT  1.780 2.310 1.800 2.640 ;
        RECT  1.800 2.310 1.880 2.630 ;
        RECT  1.880 2.310 2.980 2.550 ;
        RECT  2.980 2.310 3.380 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.160 2.820 2.630 3.250 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.450 5.440 ;
        RECT  0.450 4.000 0.460 5.440 ;
        RECT  0.460 3.800 0.860 5.440 ;
        RECT  0.860 4.000 0.870 5.440 ;
        RECT  0.870 4.640 4.090 5.440 ;
        RECT  4.090 4.210 4.100 5.440 ;
        RECT  4.100 4.010 4.500 5.440 ;
        RECT  4.500 4.210 4.510 5.440 ;
        RECT  4.510 4.640 5.360 5.440 ;
        RECT  5.360 4.210 5.370 5.440 ;
        RECT  5.370 4.010 5.770 5.440 ;
        RECT  5.770 4.210 5.780 5.440 ;
        RECT  5.780 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.050 0.400 ;
        RECT  1.050 -0.400 1.450 0.560 ;
        RECT  1.450 -0.400 2.720 0.400 ;
        RECT  2.720 -0.400 3.120 0.560 ;
        RECT  3.120 -0.400 4.080 0.400 ;
        RECT  4.080 -0.400 4.090 0.670 ;
        RECT  4.090 -0.400 4.490 0.870 ;
        RECT  4.490 -0.400 4.500 0.670 ;
        RECT  4.500 -0.400 5.360 0.400 ;
        RECT  5.360 -0.400 5.370 0.670 ;
        RECT  5.370 -0.400 5.770 0.870 ;
        RECT  5.770 -0.400 5.780 0.670 ;
        RECT  5.780 -0.400 5.940 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.220 1.150 4.460 2.240 ;
        RECT  2.270 1.150 4.220 1.390 ;
        RECT  2.260 3.700 2.660 4.100 ;
        RECT  1.870 1.110 2.270 1.510 ;
        RECT  1.820 3.700 2.260 3.940 ;
        RECT  0.570 1.110 1.870 1.350 ;
        RECT  1.580 3.180 1.820 3.940 ;
        RECT  0.410 3.180 1.580 3.420 ;
        RECT  0.410 0.940 0.570 1.350 ;
        RECT  0.170 0.940 0.410 3.420 ;
    END
END OR3X4

MACRO OR3X2
    CLASS CORE ;
    FOREIGN OR3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OR3XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.000 3.130 3.400 4.110 ;
        RECT  3.390 0.660 3.500 1.840 ;
        RECT  3.400 3.130 3.510 3.370 ;
        RECT  3.500 0.660 3.510 2.090 ;
        RECT  3.510 0.660 3.750 3.370 ;
        RECT  3.750 0.660 3.760 2.090 ;
        RECT  3.760 0.660 3.790 1.840 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.870 2.370 2.440 2.790 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.410 1.730 1.930 2.100 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.380 1.210 2.780 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 2.180 5.440 ;
        RECT  2.180 4.480 2.580 5.440 ;
        RECT  2.580 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.930 0.400 ;
        RECT  0.930 -0.400 1.330 0.560 ;
        RECT  1.330 -0.400 2.560 0.400 ;
        RECT  2.560 -0.400 2.570 0.410 ;
        RECT  2.570 -0.400 2.970 0.560 ;
        RECT  2.970 -0.400 2.980 0.410 ;
        RECT  2.980 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.820 1.060 3.060 2.310 ;
        RECT  0.400 1.060 2.820 1.460 ;
        RECT  0.400 3.070 0.750 3.470 ;
        RECT  0.170 1.060 0.400 3.470 ;
        RECT  0.160 1.070 0.170 3.470 ;
    END
END OR3X2

MACRO OR3X1
    CLASS CORE ;
    FOREIGN OR3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OR3XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.000 3.080 3.400 3.480 ;
        RECT  3.400 3.080 3.510 3.320 ;
        RECT  3.500 1.830 3.510 2.090 ;
        RECT  3.390 1.010 3.510 1.410 ;
        RECT  3.510 1.010 3.750 3.320 ;
        RECT  3.750 1.830 3.760 2.090 ;
        RECT  3.750 1.010 3.790 1.410 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.870 2.360 2.440 2.800 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.400 1.580 1.870 2.090 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.230 1.080 2.650 ;
        RECT  1.080 2.390 1.120 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 2.180 5.440 ;
        RECT  2.180 4.480 2.580 5.440 ;
        RECT  2.580 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.960 0.400 ;
        RECT  0.960 -0.400 1.360 0.560 ;
        RECT  1.360 -0.400 2.580 0.400 ;
        RECT  2.580 -0.400 2.980 0.560 ;
        RECT  2.980 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.970 1.690 3.140 2.090 ;
        RECT  2.740 1.070 2.970 2.090 ;
        RECT  2.730 1.070 2.740 2.010 ;
        RECT  2.110 1.070 2.730 1.310 ;
        RECT  1.710 0.910 2.110 1.310 ;
        RECT  0.570 1.070 1.710 1.310 ;
        RECT  0.440 2.960 0.840 3.360 ;
        RECT  0.490 0.910 0.570 1.310 ;
        RECT  0.400 0.900 0.490 1.310 ;
        RECT  0.400 2.960 0.440 3.200 ;
        RECT  0.160 0.900 0.400 3.200 ;
    END
END OR3X1

MACRO OR2XL
    CLASS CORE ;
    FOREIGN OR2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.060 3.270 2.090 3.670 ;
        RECT  2.090 3.220 2.180 3.670 ;
        RECT  2.070 1.390 2.190 1.790 ;
        RECT  2.180 2.950 2.230 3.670 ;
        RECT  2.190 1.390 2.230 1.840 ;
        RECT  2.230 1.390 2.470 3.670 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.380 1.220 3.220 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.160 1.830 0.580 2.530 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.080 5.440 ;
        RECT  1.080 4.480 1.480 5.440 ;
        RECT  1.480 4.640 2.640 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.440 0.400 ;
        RECT  0.440 -0.400 1.420 0.560 ;
        RECT  1.420 -0.400 2.640 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.780 2.120 1.930 2.520 ;
        RECT  1.540 1.270 1.780 3.810 ;
        RECT  0.460 1.270 1.540 1.510 ;
        RECT  0.570 3.570 1.540 3.810 ;
        RECT  0.170 3.490 0.570 3.890 ;
    END
END OR2XL

MACRO OR2X4
    CLASS CORE ;
    FOREIGN OR2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OR2XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.720 1.150 2.750 1.550 ;
        RECT  2.750 1.150 2.760 2.660 ;
        RECT  2.760 1.140 2.780 2.660 ;
        RECT  2.780 1.140 2.790 2.950 ;
        RECT  2.790 1.140 3.180 3.150 ;
        RECT  3.180 1.260 3.190 3.150 ;
        RECT  3.190 1.380 3.200 2.950 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.450 1.630 1.870 2.100 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.730 2.380 0.740 2.660 ;
        RECT  0.740 2.070 1.140 2.660 ;
        RECT  1.140 2.380 1.150 2.660 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 2.150 5.440 ;
        RECT  2.150 4.020 2.550 5.440 ;
        RECT  2.550 4.640 3.400 5.440 ;
        RECT  3.400 4.020 3.800 5.440 ;
        RECT  3.800 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.320 0.400 ;
        RECT  0.320 -0.400 0.740 1.550 ;
        RECT  0.740 1.140 0.780 1.540 ;
        RECT  0.740 -0.400 1.990 0.400 ;
        RECT  1.990 -0.400 2.390 0.560 ;
        RECT  2.390 -0.400 3.390 0.400 ;
        RECT  3.390 -0.400 3.790 0.560 ;
        RECT  3.790 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.460 2.070 3.700 3.670 ;
        RECT  2.380 3.430 3.460 3.670 ;
        RECT  2.140 1.030 2.380 3.670 ;
        RECT  1.580 1.030 2.140 1.270 ;
        RECT  1.210 3.320 2.140 3.670 ;
        RECT  1.180 0.890 1.580 1.290 ;
        RECT  0.810 3.020 1.210 4.000 ;
    END
END OR2X4

MACRO OR2X2
    CLASS CORE ;
    FOREIGN OR2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OR2XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 3.510 2.280 3.770 ;
        RECT  2.280 3.510 2.820 3.920 ;
        RECT  2.700 1.030 2.820 1.430 ;
        RECT  2.820 1.030 2.970 3.920 ;
        RECT  2.970 1.030 3.060 3.750 ;
        RECT  3.060 1.030 3.100 1.430 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.160 1.710 1.220 2.110 ;
        RECT  1.220 1.700 1.560 2.110 ;
        RECT  1.560 1.700 1.800 2.100 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.420 2.170 0.820 2.630 ;
        RECT  0.820 2.390 0.860 2.630 ;
        RECT  0.860 2.390 1.120 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.460 5.440 ;
        RECT  1.460 4.480 1.860 5.440 ;
        RECT  1.860 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.180 1.240 ;
        RECT  0.180 -0.400 0.580 1.440 ;
        RECT  0.580 -0.400 0.590 1.240 ;
        RECT  0.590 -0.400 1.760 0.400 ;
        RECT  1.760 -0.400 1.770 0.410 ;
        RECT  1.770 -0.400 2.170 0.560 ;
        RECT  2.170 -0.400 2.180 0.410 ;
        RECT  2.180 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.380 2.080 2.540 2.480 ;
        RECT  2.140 1.150 2.380 3.200 ;
        RECT  1.340 1.150 2.140 1.390 ;
        RECT  0.580 2.960 2.140 3.200 ;
        RECT  0.940 1.030 1.340 1.430 ;
        RECT  0.180 2.960 0.580 3.400 ;
    END
END OR2X2

MACRO OR2X1
    CLASS CORE ;
    FOREIGN OR2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OR2XL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.060 3.270 2.090 3.670 ;
        RECT  2.090 3.220 2.180 3.670 ;
        RECT  2.070 1.290 2.190 1.690 ;
        RECT  2.180 2.950 2.230 3.670 ;
        RECT  2.190 1.290 2.230 1.840 ;
        RECT  2.230 1.290 2.470 3.670 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.380 1.220 3.220 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.160 1.830 0.580 2.500 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.080 5.440 ;
        RECT  1.080 4.480 1.480 5.440 ;
        RECT  1.480 4.640 2.640 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.300 0.400 ;
        RECT  0.300 -0.400 1.280 0.560 ;
        RECT  1.280 -0.400 2.640 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.780 2.120 1.930 2.520 ;
        RECT  1.540 1.310 1.780 3.810 ;
        RECT  0.850 1.310 1.540 1.550 ;
        RECT  0.570 3.570 1.540 3.810 ;
        RECT  0.440 1.260 0.850 1.550 ;
        RECT  0.170 3.490 0.570 3.890 ;
    END
END OR2X1

MACRO OAI33XL
    CLASS CORE ;
    FOREIGN OAI33XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.260 3.490 2.970 3.890 ;
        RECT  3.130 1.460 3.140 1.920 ;
        RECT  3.140 1.250 3.410 1.920 ;
        RECT  3.410 1.250 3.540 1.910 ;
        RECT  3.540 1.670 4.660 1.910 ;
        RECT  2.970 3.490 4.830 3.730 ;
        RECT  4.820 2.390 4.830 2.650 ;
        RECT  4.660 1.120 4.830 1.910 ;
        RECT  4.830 1.120 5.070 3.730 ;
        RECT  5.070 2.390 5.080 2.650 ;
        END
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.510 3.180 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 1.120 2.650 ;
        RECT  1.120 2.390 1.190 2.630 ;
        RECT  1.190 2.220 1.430 2.630 ;
        RECT  1.430 2.220 1.590 2.620 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.940 1.900 3.220 ;
        RECT  1.900 2.650 2.300 3.220 ;
        RECT  2.300 2.940 2.310 3.220 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 2.360 4.470 3.210 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.410 2.180 3.850 2.660 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.620 2.650 2.840 3.050 ;
        RECT  2.840 2.650 3.090 3.210 ;
        RECT  3.090 2.950 3.100 3.210 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.420 5.440 ;
        RECT  0.420 4.480 0.820 5.440 ;
        RECT  0.820 4.640 4.100 5.440 ;
        RECT  4.100 4.480 4.500 5.440 ;
        RECT  4.500 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.610 0.400 ;
        RECT  1.610 -0.400 1.620 1.270 ;
        RECT  1.620 -0.400 2.020 1.390 ;
        RECT  2.020 -0.400 2.030 1.270 ;
        RECT  2.030 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.140 1.150 4.300 1.390 ;
        RECT  3.900 0.730 4.140 1.390 ;
        RECT  2.780 0.730 3.900 0.970 ;
        RECT  2.620 0.730 2.780 1.540 ;
        RECT  2.540 0.730 2.620 1.910 ;
        RECT  2.380 1.140 2.540 1.910 ;
        RECT  1.260 1.670 2.380 1.910 ;
        RECT  1.020 1.140 1.260 1.910 ;
        RECT  0.860 1.140 1.020 1.540 ;
    END
END OAI33XL

MACRO OAI33X4
    CLASS CORE ;
    FOREIGN OAI33X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI33XL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.870 2.940 5.270 3.340 ;
        RECT  5.270 2.940 5.390 3.220 ;
        RECT  5.180 1.390 5.390 1.630 ;
        RECT  5.390 1.390 5.630 3.220 ;
        RECT  5.630 1.820 5.830 3.220 ;
        END
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.630 2.550 3.790 2.950 ;
        RECT  3.790 2.550 4.030 3.180 ;
        RECT  4.030 2.940 4.160 3.180 ;
        RECT  4.160 2.940 4.400 3.210 ;
        RECT  4.400 2.950 4.420 3.210 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.310 1.820 3.500 2.220 ;
        RECT  3.500 1.810 3.870 2.230 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.470 2.460 2.630 2.860 ;
        RECT  2.630 2.460 2.840 3.200 ;
        RECT  2.840 2.460 2.870 3.210 ;
        RECT  2.870 2.950 3.100 3.210 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.670 0.460 2.090 ;
        RECT  0.460 1.670 0.690 2.080 ;
        RECT  0.690 1.680 0.810 2.080 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.380 1.280 2.660 ;
        RECT  1.280 2.020 1.520 2.660 ;
        RECT  1.520 2.380 1.530 2.660 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.460 4.060 2.290 4.370 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.410 5.440 ;
        RECT  0.410 4.480 0.810 5.440 ;
        RECT  0.810 4.640 3.940 5.440 ;
        RECT  3.940 4.480 4.340 5.440 ;
        RECT  4.340 4.640 5.600 5.440 ;
        RECT  5.600 4.210 6.000 5.440 ;
        RECT  6.000 4.640 7.260 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 2.970 0.400 ;
        RECT  2.970 -0.400 3.370 0.560 ;
        RECT  3.370 -0.400 4.490 0.400 ;
        RECT  4.490 -0.400 4.890 0.560 ;
        RECT  4.890 -0.400 5.890 0.400 ;
        RECT  5.890 -0.400 6.290 0.560 ;
        RECT  6.290 -0.400 7.260 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  7.020 0.870 7.090 1.460 ;
        RECT  6.780 0.870 7.020 3.740 ;
        RECT  6.690 0.870 6.780 1.460 ;
        RECT  4.870 0.870 6.690 1.110 ;
        RECT  6.280 2.580 6.520 3.930 ;
        RECT  3.700 3.690 6.280 3.930 ;
        RECT  4.870 2.140 5.150 2.540 ;
        RECT  4.750 0.870 4.870 2.540 ;
        RECT  4.630 0.870 4.750 2.380 ;
        RECT  3.970 1.070 4.170 1.470 ;
        RECT  2.550 1.060 3.970 1.480 ;
        RECT  3.460 3.490 3.700 3.930 ;
        RECT  2.070 3.490 3.460 3.730 ;
        RECT  2.350 1.070 2.550 1.470 ;
        RECT  1.830 1.070 2.070 3.730 ;
        RECT  1.590 1.070 1.830 1.470 ;
        RECT  0.170 1.160 1.590 1.400 ;
    END
END OAI33X4

MACRO OAI33X2
    CLASS CORE ;
    FOREIGN OAI33X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI33XL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.960 4.130 3.090 4.370 ;
        RECT  3.090 4.080 3.180 4.370 ;
        RECT  3.180 3.940 3.420 4.370 ;
        RECT  3.420 3.940 5.500 4.180 ;
        RECT  5.500 3.830 5.900 4.180 ;
        RECT  5.900 3.940 6.140 4.180 ;
        RECT  6.140 3.940 6.400 4.330 ;
        RECT  6.400 3.940 7.470 4.180 ;
        RECT  7.470 3.760 7.520 4.180 ;
        RECT  4.500 1.270 7.520 1.510 ;
        RECT  7.520 1.270 7.760 4.180 ;
        END
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.460 2.990 ;
        RECT  0.460 2.400 0.920 2.990 ;
        RECT  0.920 2.740 1.160 3.730 ;
        RECT  1.160 3.490 2.580 3.730 ;
        RECT  2.580 3.420 2.820 3.730 ;
        RECT  2.820 3.420 3.500 3.660 ;
        RECT  3.500 2.660 3.740 3.660 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.260 2.220 2.840 2.460 ;
        RECT  2.840 2.220 3.100 2.650 ;
        RECT  3.100 2.220 3.110 2.640 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.930 1.780 3.210 ;
        RECT  1.780 2.930 1.980 3.200 ;
        RECT  1.980 2.740 2.220 3.200 ;
        RECT  2.220 2.740 2.380 2.980 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.510 2.090 ;
        RECT  3.510 1.830 3.760 2.260 ;
        RECT  3.760 2.020 4.070 2.260 ;
        RECT  4.070 2.020 4.080 2.380 ;
        RECT  4.080 2.020 4.320 3.480 ;
        RECT  4.320 3.200 4.510 3.480 ;
        RECT  4.510 3.240 6.710 3.480 ;
        RECT  6.710 3.200 7.000 3.480 ;
        RECT  7.000 2.430 7.280 3.480 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.820 1.830 4.870 2.090 ;
        RECT  4.870 1.830 5.080 2.360 ;
        RECT  5.080 1.840 5.110 2.360 ;
        RECT  5.110 1.840 6.290 2.080 ;
        RECT  6.290 1.840 6.530 2.430 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.470 2.390 5.890 2.970 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.220 5.440 ;
        RECT  0.220 4.480 0.620 5.440 ;
        RECT  0.620 4.640 3.700 5.440 ;
        RECT  3.700 4.480 4.100 5.440 ;
        RECT  4.100 4.640 7.240 5.440 ;
        RECT  7.240 4.480 7.640 5.440 ;
        RECT  7.640 4.640 7.920 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.360 0.400 ;
        RECT  0.360 -0.400 0.370 0.860 ;
        RECT  0.370 -0.400 0.770 1.060 ;
        RECT  0.770 -0.400 0.780 0.860 ;
        RECT  0.780 -0.400 2.050 0.400 ;
        RECT  2.050 -0.400 2.060 0.730 ;
        RECT  2.060 -0.400 2.460 0.930 ;
        RECT  2.460 -0.400 2.470 0.730 ;
        RECT  2.470 -0.400 7.920 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.600 0.670 7.430 0.910 ;
        RECT  4.360 0.670 4.600 0.920 ;
        RECT  3.290 0.680 4.360 0.920 ;
        RECT  3.290 1.310 3.350 1.550 ;
        RECT  3.050 0.680 3.290 1.550 ;
        RECT  1.640 1.310 3.050 1.550 ;
        RECT  1.240 1.310 1.640 1.790 ;
    END
END OAI33X2

MACRO OAI33X1
    CLASS CORE ;
    FOREIGN OAI33X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI33XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.170 3.490 2.570 3.890 ;
        RECT  2.570 3.490 2.970 3.780 ;
        RECT  3.130 1.680 3.140 1.920 ;
        RECT  3.140 1.470 3.410 1.920 ;
        RECT  3.410 1.470 3.540 1.910 ;
        RECT  3.540 1.670 4.660 1.910 ;
        RECT  2.970 3.490 4.830 3.730 ;
        RECT  4.820 2.390 4.830 2.650 ;
        RECT  4.660 1.390 4.830 1.910 ;
        RECT  4.830 1.390 5.060 3.730 ;
        RECT  5.060 1.520 5.070 3.730 ;
        RECT  5.070 2.390 5.080 2.650 ;
        END
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.510 3.180 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 1.100 2.650 ;
        RECT  1.100 2.220 1.120 2.650 ;
        RECT  1.120 2.220 1.500 2.640 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.950 1.780 3.210 ;
        RECT  1.780 2.950 1.860 3.190 ;
        RECT  1.860 2.270 2.100 3.190 ;
        RECT  2.100 2.270 2.260 2.670 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 2.360 4.470 3.210 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.410 2.180 3.850 2.660 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.670 2.270 2.750 2.670 ;
        RECT  2.750 2.270 3.090 3.210 ;
        RECT  3.090 2.950 3.100 3.210 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 4.150 5.440 ;
        RECT  4.150 4.480 4.550 5.440 ;
        RECT  4.550 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.610 0.400 ;
        RECT  1.610 -0.400 1.620 1.270 ;
        RECT  1.620 -0.400 2.020 1.390 ;
        RECT  2.020 -0.400 2.030 1.270 ;
        RECT  2.030 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.900 0.940 4.300 1.390 ;
        RECT  2.780 0.940 3.900 1.180 ;
        RECT  2.620 0.940 2.780 1.540 ;
        RECT  2.380 0.940 2.620 1.910 ;
        RECT  1.260 1.670 2.380 1.910 ;
        RECT  1.020 1.140 1.260 1.910 ;
        RECT  0.860 1.140 1.020 1.540 ;
    END
END OAI33X1

MACRO OAI32XL
    CLASS CORE ;
    FOREIGN OAI32XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.050 3.490 2.450 3.890 ;
        RECT  3.200 1.460 3.210 1.920 ;
        RECT  3.210 1.250 3.510 1.920 ;
        RECT  3.510 1.250 3.610 1.910 ;
        RECT  2.450 3.490 4.170 3.730 ;
        RECT  4.160 2.390 4.170 2.650 ;
        RECT  3.610 1.670 4.170 1.910 ;
        RECT  4.170 1.670 4.410 3.730 ;
        RECT  4.410 2.390 4.420 2.650 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.450 2.390 3.780 3.050 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.950 2.850 3.210 ;
        RECT  2.690 2.200 2.850 2.600 ;
        RECT  2.850 2.200 3.090 3.210 ;
        RECT  3.090 2.950 3.100 3.210 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.510 3.180 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 1.120 2.650 ;
        RECT  1.120 2.390 1.180 2.630 ;
        RECT  1.180 2.220 1.420 2.630 ;
        RECT  1.420 2.220 1.580 2.620 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.950 1.780 3.210 ;
        RECT  1.780 2.950 1.860 3.190 ;
        RECT  1.860 2.650 2.260 3.190 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 3.340 5.440 ;
        RECT  3.340 4.480 3.740 5.440 ;
        RECT  3.740 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 1.320 ;
        RECT  0.170 -0.400 0.570 1.520 ;
        RECT  0.570 -0.400 0.580 1.320 ;
        RECT  0.580 -0.400 1.680 0.400 ;
        RECT  1.680 -0.400 1.690 1.270 ;
        RECT  1.690 -0.400 2.090 1.390 ;
        RECT  2.090 -0.400 2.100 1.270 ;
        RECT  2.100 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.220 1.150 4.380 1.390 ;
        RECT  3.980 0.730 4.220 1.390 ;
        RECT  2.850 0.730 3.980 0.970 ;
        RECT  2.690 0.730 2.850 1.540 ;
        RECT  2.610 0.730 2.690 1.910 ;
        RECT  2.450 1.140 2.610 1.910 ;
        RECT  1.330 1.670 2.450 1.910 ;
        RECT  1.090 1.120 1.330 1.910 ;
        RECT  0.930 1.120 1.090 1.520 ;
    END
END OAI32XL

MACRO OAI32X4
    CLASS CORE ;
    FOREIGN OAI32X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI32XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.210 2.940 4.730 3.340 ;
        RECT  4.470 1.390 4.730 1.630 ;
        RECT  4.730 1.390 5.160 3.340 ;
        RECT  5.160 1.390 5.170 3.220 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.460 2.980 ;
        RECT  0.460 2.400 0.630 2.980 ;
        RECT  0.630 2.620 0.640 2.980 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 3.510 1.070 3.770 ;
        RECT  1.070 3.510 1.120 4.340 ;
        RECT  1.120 3.520 1.310 4.340 ;
        RECT  1.310 3.940 1.660 4.340 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.060 2.550 3.420 2.950 ;
        RECT  3.420 2.550 3.460 3.200 ;
        RECT  3.460 2.630 3.500 3.200 ;
        RECT  3.500 2.630 3.660 3.210 ;
        RECT  3.660 2.950 3.760 3.210 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.580 1.820 2.770 2.220 ;
        RECT  2.770 1.810 3.140 2.230 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.390 1.870 2.650 ;
        RECT  1.870 2.310 2.270 2.710 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 3.360 5.440 ;
        RECT  3.360 4.480 3.760 5.440 ;
        RECT  3.760 4.640 5.020 5.440 ;
        RECT  5.020 4.210 5.420 5.440 ;
        RECT  5.420 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 2.240 0.400 ;
        RECT  2.240 -0.400 2.640 0.560 ;
        RECT  2.640 -0.400 3.800 0.400 ;
        RECT  3.800 -0.400 4.200 0.560 ;
        RECT  4.200 -0.400 5.200 0.400 ;
        RECT  5.200 -0.400 5.600 0.560 ;
        RECT  5.600 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.360 1.060 6.400 1.460 ;
        RECT  6.330 0.870 6.360 1.460 ;
        RECT  6.090 0.870 6.330 3.740 ;
        RECT  6.000 0.870 6.090 1.460 ;
        RECT  4.190 0.870 6.000 1.110 ;
        RECT  5.610 2.580 5.850 3.930 ;
        RECT  3.040 3.690 5.610 3.930 ;
        RECT  4.190 1.910 4.490 2.310 ;
        RECT  4.090 0.870 4.190 2.310 ;
        RECT  3.950 0.870 4.090 2.150 ;
        RECT  3.260 1.070 3.460 1.470 ;
        RECT  1.820 1.060 3.260 1.480 ;
        RECT  2.800 3.350 3.040 3.930 ;
        RECT  1.990 3.350 2.800 3.590 ;
        RECT  1.590 2.990 1.990 3.590 ;
        RECT  1.620 1.070 1.820 1.470 ;
        RECT  1.160 2.990 1.590 3.230 ;
        RECT  1.160 1.070 1.230 1.470 ;
        RECT  0.920 1.070 1.160 3.230 ;
        RECT  0.830 1.070 0.920 1.470 ;
    END
END OAI32X4

MACRO OAI32X2
    CLASS CORE ;
    FOREIGN OAI32X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI32XL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.960 4.130 3.090 4.370 ;
        RECT  3.090 4.080 3.100 4.370 ;
        RECT  3.100 3.940 3.340 4.370 ;
        RECT  3.340 3.940 5.220 4.180 ;
        RECT  5.220 3.600 5.620 4.180 ;
        RECT  5.620 3.940 6.050 4.180 ;
        RECT  6.050 3.510 6.380 4.180 ;
        RECT  3.900 1.470 6.380 1.710 ;
        RECT  6.380 1.470 6.620 4.180 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 2.390 4.170 2.650 ;
        RECT  4.170 1.990 4.420 2.650 ;
        RECT  4.420 1.990 4.640 2.400 ;
        RECT  4.640 1.990 5.700 2.230 ;
        RECT  5.700 1.990 6.100 2.320 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.820 2.950 4.970 3.210 ;
        RECT  4.970 2.520 5.080 3.210 ;
        RECT  5.080 2.520 5.210 3.200 ;
        RECT  5.210 2.520 5.380 2.760 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.460 2.990 ;
        RECT  0.460 2.400 0.920 2.990 ;
        RECT  0.920 2.740 1.160 3.730 ;
        RECT  1.160 3.490 2.580 3.730 ;
        RECT  2.580 3.420 2.820 3.730 ;
        RECT  2.820 3.420 3.410 3.660 ;
        RECT  3.410 3.220 3.470 3.660 ;
        RECT  3.470 2.670 3.710 3.660 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.260 2.220 2.840 2.460 ;
        RECT  2.840 2.220 3.100 2.650 ;
        RECT  3.100 2.220 3.110 2.640 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.930 1.780 3.210 ;
        RECT  1.780 2.930 1.980 3.200 ;
        RECT  1.980 2.740 2.220 3.200 ;
        RECT  2.220 2.740 2.380 2.980 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.220 5.440 ;
        RECT  0.220 4.480 0.620 5.440 ;
        RECT  0.620 4.640 3.700 5.440 ;
        RECT  3.700 4.480 4.100 5.440 ;
        RECT  4.100 4.640 6.500 5.440 ;
        RECT  6.500 4.480 6.900 5.440 ;
        RECT  6.900 4.640 7.260 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.420 0.400 ;
        RECT  0.420 -0.400 0.430 0.860 ;
        RECT  0.430 -0.400 0.830 1.060 ;
        RECT  0.830 -0.400 0.840 0.860 ;
        RECT  0.840 -0.400 2.110 0.400 ;
        RECT  2.110 -0.400 2.120 0.860 ;
        RECT  2.120 -0.400 2.520 1.060 ;
        RECT  2.520 -0.400 2.530 0.860 ;
        RECT  2.530 -0.400 7.260 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.410 0.740 5.120 0.980 ;
        RECT  3.210 0.740 3.410 1.790 ;
        RECT  3.170 0.740 3.210 1.800 ;
        RECT  1.440 1.380 3.170 1.800 ;
        RECT  1.240 1.390 1.440 1.790 ;
    END
END OAI32X2

MACRO OAI32X1
    CLASS CORE ;
    FOREIGN OAI32X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI32XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.050 3.490 2.450 3.890 ;
        RECT  3.210 1.480 3.370 1.720 ;
        RECT  3.370 1.480 3.610 1.910 ;
        RECT  2.450 3.490 4.170 3.730 ;
        RECT  4.160 2.390 4.170 2.650 ;
        RECT  3.610 1.670 4.170 1.910 ;
        RECT  4.170 1.670 4.410 3.730 ;
        RECT  4.410 2.390 4.420 2.650 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.450 2.310 3.780 2.910 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.690 2.420 2.750 2.820 ;
        RECT  2.750 2.420 3.090 3.210 ;
        RECT  3.090 2.950 3.100 3.210 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.210 2.650 ;
        RECT  0.210 2.390 0.500 3.180 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 1.120 2.650 ;
        RECT  1.120 2.390 1.140 2.630 ;
        RECT  1.140 2.220 1.540 2.630 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.950 1.780 3.210 ;
        RECT  1.780 2.950 1.860 3.190 ;
        RECT  1.860 2.650 2.260 3.190 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 3.340 5.440 ;
        RECT  3.340 4.480 3.740 5.440 ;
        RECT  3.740 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 1.420 ;
        RECT  0.170 -0.400 0.570 1.620 ;
        RECT  0.570 -0.400 0.580 1.420 ;
        RECT  0.580 -0.400 1.680 0.400 ;
        RECT  1.680 -0.400 1.690 1.270 ;
        RECT  1.690 -0.400 2.090 1.390 ;
        RECT  2.090 -0.400 2.100 1.270 ;
        RECT  2.100 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.980 0.940 4.380 1.390 ;
        RECT  2.850 0.940 3.980 1.180 ;
        RECT  2.690 0.940 2.850 1.540 ;
        RECT  2.450 0.940 2.690 1.910 ;
        RECT  1.330 1.670 2.450 1.910 ;
        RECT  1.090 1.140 1.330 1.910 ;
        RECT  0.930 1.140 1.090 1.540 ;
    END
END OAI32X1

MACRO OAI31XL
    CLASS CORE ;
    FOREIGN OAI31XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.920 3.090 2.320 3.490 ;
        RECT  3.390 1.160 3.410 1.560 ;
        RECT  3.410 1.160 3.500 1.840 ;
        RECT  2.320 3.090 3.510 3.330 ;
        RECT  3.500 1.160 3.510 2.090 ;
        RECT  3.510 1.160 3.750 3.330 ;
        RECT  3.750 1.160 3.760 2.090 ;
        RECT  3.760 1.160 3.790 1.840 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.750 2.090 3.150 2.700 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.990 0.460 2.650 ;
        RECT  0.460 1.990 0.500 2.530 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 1.120 2.090 ;
        RECT  1.120 1.840 1.630 2.080 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.390 1.540 2.650 ;
        RECT  1.540 2.380 1.780 2.650 ;
        RECT  1.780 2.380 1.950 2.620 ;
        RECT  1.950 1.850 2.190 2.620 ;
        RECT  2.190 1.850 2.350 2.250 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 2.870 5.440 ;
        RECT  2.870 4.480 3.270 5.440 ;
        RECT  3.270 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 1.800 0.400 ;
        RECT  1.800 -0.400 1.810 0.410 ;
        RECT  1.810 -0.400 2.210 0.560 ;
        RECT  2.210 -0.400 2.220 0.410 ;
        RECT  2.220 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.630 1.160 3.030 1.560 ;
        RECT  0.990 1.250 2.630 1.490 ;
    END
END OAI31XL

MACRO OAI31X4
    CLASS CORE ;
    FOREIGN OAI31X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI31XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.550 2.940 3.950 3.340 ;
        RECT  3.950 2.940 4.070 3.220 ;
        RECT  3.770 1.390 4.070 1.630 ;
        RECT  4.070 1.390 4.410 3.220 ;
        RECT  4.410 1.820 4.510 3.220 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.600 3.890 1.520 4.130 ;
        RECT  1.520 3.890 1.770 4.330 ;
        RECT  1.770 4.070 1.780 4.330 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.400 2.550 2.760 2.950 ;
        RECT  2.760 2.550 2.840 3.200 ;
        RECT  2.840 2.550 3.000 3.210 ;
        RECT  3.000 2.950 3.100 3.210 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.920 1.820 2.110 2.220 ;
        RECT  2.110 1.810 2.480 2.230 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 1.140 2.650 ;
        RECT  1.140 2.390 1.600 2.870 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 2.700 5.440 ;
        RECT  2.700 4.480 3.100 5.440 ;
        RECT  3.100 4.640 4.330 5.440 ;
        RECT  4.330 4.330 4.340 5.440 ;
        RECT  4.340 4.210 4.740 5.440 ;
        RECT  4.740 4.330 4.750 5.440 ;
        RECT  4.750 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.690 0.400 ;
        RECT  1.690 -0.400 2.090 0.560 ;
        RECT  2.090 -0.400 3.040 0.400 ;
        RECT  3.040 -0.400 3.440 0.560 ;
        RECT  3.440 -0.400 4.480 0.400 ;
        RECT  4.480 -0.400 4.880 0.560 ;
        RECT  4.880 -0.400 5.940 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.580 0.870 5.700 1.460 ;
        RECT  5.340 0.870 5.580 3.740 ;
        RECT  5.300 0.870 5.340 1.460 ;
        RECT  3.480 0.870 5.300 1.110 ;
        RECT  4.810 2.350 5.050 3.930 ;
        RECT  2.380 3.690 4.810 3.930 ;
        RECT  3.480 1.910 3.800 2.310 ;
        RECT  3.240 0.870 3.480 2.310 ;
        RECT  2.580 1.070 2.780 1.470 ;
        RECT  1.130 1.060 2.580 1.480 ;
        RECT  2.140 3.270 2.380 3.930 ;
        RECT  0.500 3.270 2.140 3.510 ;
        RECT  0.930 1.070 1.130 1.470 ;
        RECT  0.500 1.070 0.570 1.470 ;
        RECT  0.260 1.070 0.500 3.510 ;
        RECT  0.170 1.070 0.260 1.470 ;
    END
END OAI31X4

MACRO OAI31X2
    CLASS CORE ;
    FOREIGN OAI31X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI31XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.970 3.450 2.370 3.850 ;
        RECT  2.370 3.530 4.410 3.770 ;
        RECT  4.410 3.500 4.510 3.770 ;
        RECT  4.510 3.500 4.530 3.780 ;
        RECT  4.530 3.450 4.780 3.850 ;
        RECT  4.780 1.870 4.930 3.850 ;
        RECT  4.930 1.870 5.020 3.770 ;
        RECT  5.020 3.480 5.070 3.770 ;
        RECT  5.020 1.870 5.070 2.110 ;
        RECT  5.070 3.510 5.080 3.770 ;
        RECT  5.070 1.820 5.230 2.110 ;
        RECT  5.230 1.360 5.470 2.110 ;
        RECT  5.470 1.360 5.630 1.600 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.310 2.380 5.830 2.800 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.410 2.400 0.550 2.640 ;
        RECT  0.550 2.400 0.570 2.660 ;
        RECT  0.570 2.400 0.810 3.170 ;
        RECT  0.810 2.930 3.940 3.170 ;
        RECT  3.940 2.410 4.100 3.170 ;
        RECT  4.100 2.400 4.160 3.170 ;
        RECT  4.160 2.390 4.180 3.170 ;
        RECT  4.180 2.390 4.420 2.650 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 0.870 2.090 ;
        RECT  0.870 1.830 1.120 2.110 ;
        RECT  1.120 1.850 1.530 2.110 ;
        RECT  1.530 1.870 3.120 2.110 ;
        RECT  3.120 1.870 3.520 2.210 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.840 2.380 2.530 2.660 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.230 5.440 ;
        RECT  0.230 4.480 0.630 5.440 ;
        RECT  0.630 4.640 3.710 5.440 ;
        RECT  3.710 4.480 4.110 5.440 ;
        RECT  4.110 4.640 5.440 5.440 ;
        RECT  5.440 3.780 5.680 5.440 ;
        RECT  5.680 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.770 0.400 ;
        RECT  0.770 -0.400 0.780 0.690 ;
        RECT  0.780 -0.400 1.180 0.890 ;
        RECT  1.180 -0.400 1.190 0.690 ;
        RECT  1.190 -0.400 2.090 0.400 ;
        RECT  2.090 -0.400 2.100 0.690 ;
        RECT  2.100 -0.400 2.500 0.890 ;
        RECT  2.500 -0.400 2.510 0.690 ;
        RECT  2.510 -0.400 3.700 0.400 ;
        RECT  3.700 -0.400 4.100 0.560 ;
        RECT  4.100 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.230 1.220 6.390 1.620 ;
        RECT  5.990 0.830 6.230 1.620 ;
        RECT  4.910 0.830 5.990 1.070 ;
        RECT  4.670 0.830 4.910 1.570 ;
        RECT  4.510 1.170 4.670 1.570 ;
        RECT  3.300 1.250 4.510 1.490 ;
        RECT  2.900 1.170 3.300 1.570 ;
        RECT  0.570 1.250 2.900 1.490 ;
        RECT  0.170 1.170 0.570 1.570 ;
    END
END OAI31X2

MACRO OAI31X1
    CLASS CORE ;
    FOREIGN OAI31X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI31XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.990 3.090 2.390 3.490 ;
        RECT  3.390 1.200 3.500 1.860 ;
        RECT  2.390 3.090 3.510 3.330 ;
        RECT  3.500 1.200 3.510 2.090 ;
        RECT  3.510 1.200 3.750 3.330 ;
        RECT  3.750 1.200 3.760 2.090 ;
        RECT  3.760 1.200 3.790 1.860 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.390 2.890 2.650 ;
        RECT  2.890 1.960 3.150 2.700 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.000 0.500 2.650 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 1.120 2.090 ;
        RECT  1.120 1.840 1.640 2.080 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.390 1.540 2.650 ;
        RECT  1.540 2.380 1.780 2.650 ;
        RECT  1.780 2.380 1.940 2.620 ;
        RECT  1.940 1.850 2.180 2.620 ;
        RECT  2.180 1.850 2.340 2.250 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 3.040 5.440 ;
        RECT  3.040 4.480 3.440 5.440 ;
        RECT  3.440 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 1.800 0.400 ;
        RECT  1.800 -0.400 1.810 0.410 ;
        RECT  1.810 -0.400 2.210 0.560 ;
        RECT  2.210 -0.400 2.220 0.410 ;
        RECT  2.220 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.630 1.160 3.030 1.560 ;
        RECT  0.990 1.250 2.630 1.490 ;
    END
END OAI31X1

MACRO OAI2BB2XL
    CLASS CORE ;
    FOREIGN OAI2BB2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.870 3.630 3.270 4.030 ;
        RECT  3.270 3.630 4.170 3.870 ;
        RECT  4.160 1.830 4.170 2.090 ;
        RECT  4.050 0.710 4.170 1.300 ;
        RECT  4.170 0.710 4.410 3.870 ;
        RECT  4.410 1.830 4.420 2.090 ;
        RECT  4.410 0.710 4.450 1.300 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.040 1.820 2.530 2.230 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.800 2.010 2.840 2.410 ;
        RECT  2.840 2.010 3.100 2.650 ;
        RECT  3.100 2.010 3.200 2.410 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.380 1.210 2.960 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.210 2.090 ;
        RECT  0.210 1.800 0.510 2.420 ;
        END
    END A0N
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.480 5.440 ;
        RECT  0.480 4.480 0.880 5.440 ;
        RECT  0.880 4.640 1.590 5.440 ;
        RECT  1.590 4.480 1.990 5.440 ;
        RECT  1.990 4.640 3.690 5.440 ;
        RECT  3.690 4.480 4.090 5.440 ;
        RECT  4.090 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 2.520 0.400 ;
        RECT  2.520 -0.400 2.530 0.860 ;
        RECT  2.530 -0.400 2.930 0.980 ;
        RECT  2.930 -0.400 2.940 0.860 ;
        RECT  2.940 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.560 2.740 3.800 3.350 ;
        RECT  3.530 0.720 3.690 1.120 ;
        RECT  1.720 3.110 3.560 3.350 ;
        RECT  3.290 0.720 3.530 1.550 ;
        RECT  2.250 1.310 3.290 1.550 ;
        RECT  2.010 0.740 2.250 1.550 ;
        RECT  1.770 0.740 2.010 0.980 ;
        RECT  1.480 1.400 1.720 3.730 ;
        RECT  1.290 1.400 1.480 1.800 ;
        RECT  0.490 3.490 1.480 3.730 ;
    END
END OAI2BB2XL

MACRO OAI2BB2X4
    CLASS CORE ;
    FOREIGN OAI2BB2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI2BB2XL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  5.470 0.860 8.360 1.100 ;
        RECT  8.360 0.780 8.600 1.100 ;
        RECT  4.920 3.600 9.660 3.840 ;
        RECT  9.660 3.500 10.010 3.840 ;
        RECT  8.600 0.780 10.020 1.020 ;
        RECT  10.010 2.380 10.230 3.840 ;
        RECT  10.020 0.780 10.230 1.590 ;
        RECT  10.230 0.780 10.350 3.840 ;
        RECT  10.350 0.780 10.450 3.780 ;
        RECT  10.450 0.780 10.470 2.630 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.400 2.270 3.480 2.510 ;
        RECT  3.480 2.270 3.500 2.640 ;
        RECT  3.500 2.270 3.560 2.650 ;
        RECT  3.560 2.270 3.800 2.710 ;
        RECT  3.800 2.470 8.350 2.710 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 1.830 4.170 2.090 ;
        RECT  4.170 1.830 4.420 2.160 ;
        RECT  4.420 1.920 4.630 2.160 ;
        RECT  4.630 1.920 4.870 2.190 ;
        RECT  4.870 1.950 6.730 2.190 ;
        RECT  6.730 1.940 6.970 2.190 ;
        RECT  6.970 1.940 8.910 2.180 ;
        RECT  8.910 1.940 9.150 2.380 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 1.210 2.650 ;
        RECT  1.210 2.280 1.450 2.680 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.210 2.650 ;
        RECT  0.210 1.710 0.450 2.650 ;
        RECT  0.450 2.390 0.460 2.650 ;
        RECT  0.450 1.710 0.640 2.110 ;
        RECT  0.640 1.710 0.850 1.950 ;
        RECT  0.850 0.680 1.090 1.950 ;
        RECT  1.090 0.680 2.150 0.920 ;
        RECT  2.150 0.680 2.250 1.360 ;
        RECT  2.250 0.680 2.350 2.100 ;
        RECT  2.350 0.680 2.390 2.250 ;
        RECT  2.390 0.800 2.490 2.250 ;
        RECT  2.490 1.850 2.750 2.250 ;
        END
    END A0N
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.690 0.170 5.440 ;
        RECT  0.170 3.490 0.570 5.440 ;
        RECT  0.570 3.690 0.580 5.440 ;
        RECT  0.580 4.640 1.640 5.440 ;
        RECT  1.640 4.480 2.040 5.440 ;
        RECT  2.040 4.640 2.900 5.440 ;
        RECT  2.900 4.480 4.040 5.440 ;
        RECT  4.040 4.640 5.850 5.440 ;
        RECT  5.850 4.480 6.250 5.440 ;
        RECT  6.250 4.640 7.880 5.440 ;
        RECT  7.880 4.320 7.890 5.440 ;
        RECT  7.890 4.120 8.290 5.440 ;
        RECT  8.290 4.320 8.300 5.440 ;
        RECT  8.300 4.640 9.930 5.440 ;
        RECT  9.930 4.480 10.330 5.440 ;
        RECT  10.330 4.640 11.220 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 1.060 ;
        RECT  0.170 -0.400 0.570 1.180 ;
        RECT  0.570 -0.400 0.580 1.060 ;
        RECT  0.580 -0.400 2.670 0.400 ;
        RECT  2.670 -0.400 3.070 0.560 ;
        RECT  3.070 -0.400 3.940 0.400 ;
        RECT  3.940 -0.400 3.950 0.870 ;
        RECT  3.950 -0.400 4.350 0.990 ;
        RECT  4.350 -0.400 4.360 0.870 ;
        RECT  4.360 -0.400 7.050 0.400 ;
        RECT  7.050 -0.400 7.450 0.560 ;
        RECT  7.450 -0.400 11.220 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  9.740 1.870 9.950 2.110 ;
        RECT  9.500 1.870 9.740 3.230 ;
        RECT  9.220 1.300 9.710 1.540 ;
        RECT  4.630 2.990 9.500 3.230 ;
        RECT  8.980 1.300 9.220 1.620 ;
        RECT  8.190 1.380 8.980 1.620 ;
        RECT  7.870 1.380 8.190 1.630 ;
        RECT  5.110 1.390 7.870 1.630 ;
        RECT  4.870 1.310 5.110 1.630 ;
        RECT  3.190 1.310 4.870 1.550 ;
        RECT  4.390 2.990 4.630 3.450 ;
        RECT  1.970 3.210 4.390 3.450 ;
        RECT  1.790 1.650 1.970 3.450 ;
        RECT  1.730 1.210 1.790 3.450 ;
        RECT  1.550 1.210 1.730 1.890 ;
        RECT  0.910 3.210 1.730 3.450 ;
        RECT  1.390 1.210 1.550 1.450 ;
    END
END OAI2BB2X4

MACRO OAI2BB2X2
    CLASS CORE ;
    FOREIGN OAI2BB2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI2BB2XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.910 3.940 3.310 4.340 ;
        RECT  3.310 3.940 4.550 4.180 ;
        RECT  4.370 1.300 4.830 1.700 ;
        RECT  4.550 3.940 4.950 4.340 ;
        RECT  4.950 3.940 6.050 4.180 ;
        RECT  4.830 1.460 6.050 1.700 ;
        RECT  6.050 1.460 6.140 1.860 ;
        RECT  6.050 3.780 6.150 4.180 ;
        RECT  6.140 1.460 6.150 2.090 ;
        RECT  6.150 1.460 6.390 4.180 ;
        RECT  6.390 1.830 6.400 2.090 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.250 2.390 2.490 2.920 ;
        RECT  2.490 2.680 4.150 2.920 ;
        RECT  4.150 2.680 4.390 3.660 ;
        RECT  4.390 3.420 5.390 3.660 ;
        RECT  5.390 2.970 5.480 3.660 ;
        RECT  5.480 2.950 5.540 3.660 ;
        RECT  5.540 2.390 5.630 3.660 ;
        RECT  5.630 2.390 5.780 3.210 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.820 2.200 5.080 3.100 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 0.870 2.650 ;
        RECT  0.870 2.390 1.120 2.870 ;
        RECT  1.120 2.630 1.210 2.870 ;
        RECT  1.210 2.630 1.450 3.030 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.500 2.620 ;
        END
    END A0N
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.740 0.170 5.440 ;
        RECT  0.170 3.540 0.570 5.440 ;
        RECT  0.570 3.740 0.580 5.440 ;
        RECT  0.580 4.640 1.680 5.440 ;
        RECT  1.680 3.960 1.690 5.440 ;
        RECT  1.690 3.840 2.090 5.440 ;
        RECT  2.090 3.960 2.100 5.440 ;
        RECT  2.100 4.640 3.730 5.440 ;
        RECT  3.730 4.480 4.130 5.440 ;
        RECT  4.130 4.640 5.950 5.440 ;
        RECT  5.950 4.480 6.350 5.440 ;
        RECT  6.350 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 1.190 ;
        RECT  0.170 -0.400 0.570 1.390 ;
        RECT  0.570 -0.400 0.580 1.190 ;
        RECT  0.580 -0.400 2.780 0.400 ;
        RECT  2.780 -0.400 2.790 1.110 ;
        RECT  2.790 -0.400 3.190 1.310 ;
        RECT  3.190 -0.400 3.200 1.110 ;
        RECT  3.200 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.850 1.170 4.010 1.570 ;
        RECT  3.790 3.200 3.870 3.440 ;
        RECT  3.610 1.170 3.850 1.830 ;
        RECT  3.470 3.200 3.790 3.550 ;
        RECT  2.290 1.590 3.610 1.830 ;
        RECT  1.970 3.310 3.470 3.550 ;
        RECT  2.050 1.330 2.290 1.830 ;
        RECT  1.770 2.110 1.970 3.550 ;
        RECT  1.770 0.670 1.850 0.910 ;
        RECT  1.730 0.670 1.770 3.550 ;
        RECT  1.530 0.670 1.730 2.350 ;
        RECT  1.330 3.310 1.730 3.550 ;
        RECT  1.450 0.670 1.530 0.910 ;
        RECT  1.010 3.310 1.330 3.810 ;
        RECT  0.930 3.410 1.010 3.810 ;
    END
END OAI2BB2X2

MACRO OAI2BB2X1
    CLASS CORE ;
    FOREIGN OAI2BB2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI2BB2XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.870 3.630 3.270 4.030 ;
        RECT  3.270 3.630 4.170 3.870 ;
        RECT  4.160 1.830 4.170 2.090 ;
        RECT  4.050 0.830 4.170 1.300 ;
        RECT  4.170 0.830 4.410 3.870 ;
        RECT  4.410 1.830 4.420 2.090 ;
        RECT  4.410 0.830 4.450 1.300 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.090 1.820 2.490 2.610 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.780 1.890 2.840 2.520 ;
        RECT  2.840 1.890 3.100 2.650 ;
        RECT  3.100 1.890 3.180 2.390 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.850 2.390 1.190 3.020 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.150 1.710 0.500 2.620 ;
        RECT  0.500 1.710 0.570 2.110 ;
        END
    END A0N
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.550 5.440 ;
        RECT  0.550 4.480 0.950 5.440 ;
        RECT  0.950 4.640 1.590 5.440 ;
        RECT  1.590 4.480 1.990 5.440 ;
        RECT  1.990 4.640 3.690 5.440 ;
        RECT  3.690 4.480 4.090 5.440 ;
        RECT  4.090 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 2.520 0.400 ;
        RECT  2.520 -0.400 2.530 0.860 ;
        RECT  2.530 -0.400 2.930 0.980 ;
        RECT  2.930 -0.400 2.940 0.860 ;
        RECT  2.940 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.560 2.740 3.800 3.350 ;
        RECT  3.530 0.830 3.690 1.230 ;
        RECT  1.720 3.110 3.560 3.350 ;
        RECT  3.290 0.830 3.530 1.550 ;
        RECT  2.250 1.310 3.290 1.550 ;
        RECT  2.010 0.640 2.250 1.550 ;
        RECT  1.790 0.640 2.010 0.880 ;
        RECT  1.480 1.570 1.720 3.730 ;
        RECT  1.280 1.570 1.480 1.970 ;
        RECT  0.510 3.490 1.480 3.730 ;
    END
END OAI2BB2X1

MACRO OAI2BB1XL
    CLASS CORE ;
    FOREIGN OAI2BB1XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.100 3.520 2.180 3.760 ;
        RECT  2.180 3.510 2.440 3.770 ;
        RECT  2.440 3.520 2.900 3.760 ;
        RECT  2.730 0.790 2.900 1.030 ;
        RECT  2.900 0.790 3.140 3.760 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 2.310 1.980 2.710 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.380 0.500 3.040 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.840 1.820 1.160 2.600 ;
        END
    END A0N
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 1.700 5.440 ;
        RECT  1.700 4.640 2.730 5.440 ;
        RECT  2.730 4.480 3.130 5.440 ;
        RECT  3.130 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.500 0.400 ;
        RECT  1.500 -0.400 1.510 0.910 ;
        RECT  1.510 -0.400 1.910 1.030 ;
        RECT  1.910 -0.400 1.920 0.910 ;
        RECT  1.920 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.380 1.310 2.620 3.230 ;
        RECT  0.570 1.310 2.380 1.550 ;
        RECT  1.670 2.990 2.380 3.230 ;
        RECT  1.430 2.990 1.670 3.730 ;
        RECT  0.460 3.490 1.430 3.730 ;
        RECT  0.330 0.870 0.570 1.550 ;
        RECT  0.170 0.870 0.330 1.270 ;
    END
END OAI2BB1XL

MACRO OAI2BB1X4
    CLASS CORE ;
    FOREIGN OAI2BB1X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI2BB1XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.340 2.920 3.460 3.320 ;
        RECT  3.460 2.910 4.730 3.330 ;
        RECT  2.740 0.980 4.730 1.380 ;
        RECT  4.730 0.980 4.940 3.330 ;
        RECT  4.940 0.980 5.140 3.320 ;
        RECT  5.140 0.980 5.170 3.220 ;
        RECT  5.170 0.980 5.610 1.540 ;
        RECT  5.610 0.980 5.710 1.380 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.030 2.460 2.100 2.860 ;
        RECT  2.100 1.830 2.280 2.860 ;
        RECT  2.280 1.760 2.520 2.860 ;
        RECT  2.520 1.760 3.620 2.000 ;
        RECT  3.620 1.760 3.960 2.100 ;
        RECT  3.960 1.760 4.290 2.430 ;
        RECT  4.290 2.030 4.360 2.430 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.070 0.590 2.650 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.390 1.280 1.520 2.440 ;
        RECT  1.520 1.270 1.630 2.440 ;
        RECT  1.630 1.270 1.780 1.530 ;
        END
    END A0N
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.260 0.170 5.440 ;
        RECT  0.170 4.060 0.570 5.440 ;
        RECT  0.570 4.260 0.580 5.440 ;
        RECT  0.580 4.640 1.850 5.440 ;
        RECT  1.580 3.750 1.850 4.150 ;
        RECT  1.850 3.750 2.270 5.440 ;
        RECT  2.270 3.750 2.540 4.150 ;
        RECT  2.270 4.640 3.980 5.440 ;
        RECT  3.980 4.330 3.990 5.440 ;
        RECT  3.990 4.130 4.390 5.440 ;
        RECT  4.390 4.330 4.400 5.440 ;
        RECT  4.400 4.640 5.360 5.440 ;
        RECT  5.360 4.330 5.370 5.440 ;
        RECT  5.370 4.130 5.770 5.440 ;
        RECT  5.770 4.330 5.780 5.440 ;
        RECT  5.780 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.460 0.400 ;
        RECT  1.460 -0.400 1.860 0.560 ;
        RECT  1.860 -0.400 4.020 0.400 ;
        RECT  4.020 -0.400 4.420 0.560 ;
        RECT  4.420 -0.400 5.940 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.440 2.280 5.680 3.850 ;
        RECT  3.060 3.610 5.440 3.850 ;
        RECT  3.060 2.280 3.160 2.680 ;
        RECT  2.820 2.280 3.060 3.850 ;
        RECT  1.100 3.210 2.820 3.450 ;
        RECT  0.860 1.550 1.100 3.450 ;
        RECT  0.730 1.550 0.860 1.790 ;
        RECT  0.330 1.390 0.730 1.790 ;
    END
END OAI2BB1X4

MACRO OAI2BB1X2
    CLASS CORE ;
    FOREIGN OAI2BB1X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI2BB1XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.740 1.080 2.800 1.480 ;
        RECT  2.800 1.080 3.140 1.720 ;
        RECT  3.280 2.890 3.410 3.290 ;
        RECT  3.140 1.480 3.410 1.720 ;
        RECT  3.410 2.660 3.510 3.290 ;
        RECT  3.510 2.640 3.660 3.290 ;
        RECT  3.410 1.480 3.660 1.840 ;
        RECT  3.660 1.480 3.680 3.290 ;
        RECT  3.680 1.480 3.760 3.210 ;
        RECT  3.760 1.480 3.900 3.200 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.090 1.840 2.180 2.680 ;
        RECT  2.180 1.830 2.330 2.680 ;
        RECT  2.330 1.830 2.440 2.090 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.820 0.580 2.620 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.400 1.280 1.520 2.220 ;
        RECT  1.520 1.270 1.640 2.220 ;
        RECT  1.640 1.270 1.780 1.530 ;
        END
    END A0N
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.260 5.440 ;
        RECT  0.260 4.480 0.660 5.440 ;
        RECT  0.660 4.640 2.270 5.440 ;
        RECT  2.270 4.070 2.280 5.440 ;
        RECT  2.280 3.580 2.680 5.440 ;
        RECT  2.680 4.070 2.690 5.440 ;
        RECT  2.690 4.640 3.880 5.440 ;
        RECT  3.880 4.330 3.890 5.440 ;
        RECT  3.890 4.130 4.290 5.440 ;
        RECT  4.290 4.330 4.300 5.440 ;
        RECT  4.300 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.460 0.400 ;
        RECT  1.460 -0.400 1.860 0.560 ;
        RECT  1.860 -0.400 4.020 0.400 ;
        RECT  4.020 -0.400 4.420 1.200 ;
        RECT  4.420 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.090 2.000 3.170 2.400 ;
        RECT  2.940 2.000 3.090 2.610 ;
        RECT  2.770 2.000 2.940 3.200 ;
        RECT  2.700 2.370 2.770 3.200 ;
        RECT  1.480 2.960 2.700 3.200 ;
        RECT  1.110 2.960 1.480 3.490 ;
        RECT  0.870 1.310 1.110 3.490 ;
        RECT  0.570 1.310 0.870 1.550 ;
        RECT  0.170 1.150 0.570 1.550 ;
    END
END OAI2BB1X2

MACRO OAI2BB1X1
    CLASS CORE ;
    FOREIGN OAI2BB1X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI2BB1XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.730 0.790 2.750 1.030 ;
        RECT  2.100 3.520 2.850 3.760 ;
        RECT  2.840 2.390 2.850 2.650 ;
        RECT  2.750 0.790 2.850 1.260 ;
        RECT  2.850 2.390 2.900 3.770 ;
        RECT  2.850 0.790 2.900 1.280 ;
        RECT  2.900 0.790 3.140 3.770 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.510 1.980 1.910 2.710 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.170 2.630 0.200 3.030 ;
        RECT  0.200 2.390 0.460 3.030 ;
        RECT  0.460 2.400 0.490 3.030 ;
        RECT  0.490 2.630 0.570 3.030 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.820 1.820 1.160 2.520 ;
        END
    END A0N
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 1.700 5.440 ;
        RECT  1.700 4.640 2.730 5.440 ;
        RECT  2.730 4.480 3.130 5.440 ;
        RECT  3.130 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.500 0.400 ;
        RECT  1.500 -0.400 1.510 0.910 ;
        RECT  1.510 -0.400 1.910 1.030 ;
        RECT  1.910 -0.400 1.920 0.910 ;
        RECT  1.920 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.270 1.310 2.510 3.230 ;
        RECT  0.570 1.310 2.270 1.550 ;
        RECT  1.670 2.990 2.270 3.230 ;
        RECT  1.430 2.990 1.670 3.730 ;
        RECT  0.460 3.490 1.430 3.730 ;
        RECT  0.330 0.870 0.570 1.550 ;
        RECT  0.170 0.870 0.330 1.270 ;
    END
END OAI2BB1X1

MACRO OAI22XL
    CLASS CORE ;
    FOREIGN OAI22XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.450 3.490 1.850 3.890 ;
        RECT  2.510 1.320 2.670 1.560 ;
        RECT  2.670 1.320 2.910 1.980 ;
        RECT  1.850 3.490 3.510 3.730 ;
        RECT  3.500 2.950 3.510 3.210 ;
        RECT  2.910 1.740 3.510 1.980 ;
        RECT  3.510 1.740 3.750 3.730 ;
        RECT  3.750 2.950 3.760 3.210 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.500 2.430 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 0.970 2.650 ;
        RECT  0.970 1.980 1.120 2.650 ;
        RECT  1.120 1.980 1.190 2.630 ;
        RECT  1.190 1.820 1.210 2.630 ;
        RECT  1.210 1.820 1.590 2.220 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.560 2.350 3.150 2.650 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.690 2.540 2.090 3.190 ;
        RECT  2.090 2.950 2.180 3.190 ;
        RECT  2.180 2.950 2.440 3.210 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 2.730 5.440 ;
        RECT  2.730 4.480 3.130 5.440 ;
        RECT  3.130 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.960 0.400 ;
        RECT  0.960 -0.400 1.360 0.560 ;
        RECT  1.360 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.510 1.220 3.670 1.460 ;
        RECT  3.270 0.800 3.510 1.460 ;
        RECT  2.150 0.800 3.270 1.040 ;
        RECT  1.910 0.800 2.150 1.540 ;
        RECT  1.750 1.140 1.910 1.540 ;
        RECT  0.570 1.220 1.750 1.460 ;
        RECT  0.170 1.140 0.570 1.540 ;
    END
END OAI22XL

MACRO OAI22X4
    CLASS CORE ;
    FOREIGN OAI22X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI22XL ;
    SIZE 9.900 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.300 2.940 0.700 4.050 ;
        RECT  0.700 2.940 0.980 3.220 ;
        RECT  0.980 2.940 2.880 3.180 ;
        RECT  2.880 2.940 3.280 3.920 ;
        RECT  3.280 2.940 3.650 3.220 ;
        RECT  5.100 1.220 5.300 1.620 ;
        RECT  3.650 2.940 5.580 3.180 ;
        RECT  5.580 2.940 5.980 3.920 ;
        RECT  5.980 2.940 6.280 3.230 ;
        RECT  5.300 1.210 7.880 1.630 ;
        RECT  7.880 1.210 8.090 1.920 ;
        RECT  6.280 2.940 8.180 3.180 ;
        RECT  8.090 1.220 8.290 1.920 ;
        RECT  8.290 1.420 8.300 1.920 ;
        RECT  8.180 2.940 8.580 3.920 ;
        RECT  8.580 2.940 8.690 3.340 ;
        RECT  8.300 1.500 8.690 1.920 ;
        RECT  8.690 1.500 9.130 3.340 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.920 2.420 2.980 2.660 ;
        RECT  2.980 2.380 3.860 2.660 ;
        RECT  3.860 2.190 4.260 2.660 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.560 1.900 0.860 2.300 ;
        RECT  0.860 1.830 1.120 2.300 ;
        RECT  1.120 1.900 1.200 2.300 ;
        RECT  1.200 1.900 3.140 2.140 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.610 2.070 4.620 2.660 ;
        RECT  4.620 1.900 5.170 2.660 ;
        RECT  5.170 1.900 7.110 2.140 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.840 2.420 7.460 2.660 ;
        RECT  7.460 2.380 7.700 2.660 ;
        RECT  7.700 2.380 7.720 2.650 ;
        RECT  7.720 2.380 7.940 2.620 ;
        RECT  7.940 2.190 8.180 2.620 ;
        RECT  8.180 2.190 8.340 2.590 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.570 5.440 ;
        RECT  1.570 3.970 1.580 5.440 ;
        RECT  1.580 3.480 1.980 5.440 ;
        RECT  1.980 3.970 1.990 5.440 ;
        RECT  1.990 4.640 4.240 5.440 ;
        RECT  4.240 3.970 4.250 5.440 ;
        RECT  4.250 3.480 4.650 5.440 ;
        RECT  4.650 3.970 4.660 5.440 ;
        RECT  4.660 4.640 6.850 5.440 ;
        RECT  6.850 3.970 6.860 5.440 ;
        RECT  6.860 3.480 7.260 5.440 ;
        RECT  7.260 3.970 7.270 5.440 ;
        RECT  7.270 4.640 9.900 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.830 0.400 ;
        RECT  0.830 -0.400 1.230 0.560 ;
        RECT  1.230 -0.400 2.230 0.400 ;
        RECT  2.230 -0.400 2.630 0.560 ;
        RECT  2.630 -0.400 3.630 0.400 ;
        RECT  3.630 -0.400 4.030 0.560 ;
        RECT  4.030 -0.400 9.900 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  8.840 0.990 9.040 1.230 ;
        RECT  8.600 0.680 8.840 1.230 ;
        RECT  4.710 0.680 8.600 0.920 ;
        RECT  4.470 0.680 4.710 1.620 ;
        RECT  4.310 1.220 4.470 1.620 ;
        RECT  3.310 1.300 4.310 1.540 ;
        RECT  2.910 1.220 3.310 1.620 ;
        RECT  1.910 1.300 2.910 1.540 ;
        RECT  1.510 1.220 1.910 1.620 ;
        RECT  0.490 1.220 1.510 1.460 ;
        RECT  0.250 1.220 0.490 1.620 ;
    END
END OAI22X4

MACRO OAI22X2
    CLASS CORE ;
    FOREIGN OAI22X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI22XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.170 3.610 0.570 4.010 ;
        RECT  0.570 3.610 2.430 3.850 ;
        RECT  2.430 3.520 2.530 3.850 ;
        RECT  2.530 3.500 2.750 3.850 ;
        RECT  2.750 3.500 2.760 4.060 ;
        RECT  2.760 3.120 3.160 4.100 ;
        RECT  3.160 3.610 3.510 4.100 ;
        RECT  3.780 1.210 3.960 1.610 ;
        RECT  3.960 1.210 4.200 1.850 ;
        RECT  4.200 1.610 5.300 1.850 ;
        RECT  3.510 3.610 5.520 3.850 ;
        RECT  5.300 1.210 5.700 1.850 ;
        RECT  5.700 1.520 5.830 1.850 ;
        RECT  5.520 3.610 6.150 4.020 ;
        RECT  6.140 2.390 6.150 2.650 ;
        RECT  5.830 1.610 6.150 1.850 ;
        RECT  6.150 1.610 6.390 4.020 ;
        RECT  6.390 3.630 6.400 4.020 ;
        RECT  6.390 2.390 6.400 2.650 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.180 2.390 2.160 2.790 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.210 2.090 ;
        RECT  0.210 1.830 0.430 2.110 ;
        RECT  0.430 1.830 0.460 2.430 ;
        RECT  0.460 1.870 0.830 2.430 ;
        RECT  0.830 1.870 2.560 2.110 ;
        RECT  2.560 1.870 2.960 2.470 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 2.950 4.310 3.210 ;
        RECT  4.310 2.720 4.420 3.210 ;
        RECT  4.420 2.720 4.710 3.200 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.270 2.040 3.500 2.440 ;
        RECT  3.500 2.040 3.670 2.650 ;
        RECT  3.670 2.140 3.760 2.650 ;
        RECT  3.760 2.140 5.380 2.380 ;
        RECT  5.380 2.140 5.620 2.810 ;
        RECT  5.620 2.410 5.780 2.810 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.460 5.440 ;
        RECT  1.460 4.480 1.860 5.440 ;
        RECT  1.860 4.640 4.140 5.440 ;
        RECT  4.140 4.480 4.540 5.440 ;
        RECT  4.540 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        RECT  0.980 -0.400 1.380 0.560 ;
        RECT  1.380 -0.400 2.310 0.400 ;
        RECT  2.310 -0.400 2.710 0.560 ;
        RECT  2.710 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.780 1.090 4.940 1.330 ;
        RECT  4.540 0.690 4.780 1.330 ;
        RECT  3.440 0.690 4.540 0.930 ;
        RECT  3.200 0.690 3.440 1.590 ;
        RECT  3.040 1.190 3.200 1.590 ;
        RECT  1.970 1.190 3.040 1.430 ;
        RECT  1.570 1.190 1.970 1.590 ;
        RECT  0.570 1.190 1.570 1.430 ;
        RECT  0.170 1.150 0.570 1.550 ;
    END
END OAI22X2

MACRO OAI22X1
    CLASS CORE ;
    FOREIGN OAI22X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI22XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.470 3.490 1.870 3.890 ;
        RECT  1.870 3.490 2.090 3.780 ;
        RECT  2.090 3.490 2.190 3.760 ;
        RECT  2.570 1.330 2.730 1.570 ;
        RECT  2.730 1.330 2.970 1.980 ;
        RECT  2.190 3.490 3.510 3.730 ;
        RECT  3.500 2.950 3.510 3.210 ;
        RECT  2.970 1.740 3.510 1.980 ;
        RECT  3.510 1.740 3.750 3.730 ;
        RECT  3.750 2.950 3.760 3.210 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.820 0.500 2.430 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 0.960 2.650 ;
        RECT  0.960 1.820 1.200 2.650 ;
        RECT  1.200 1.820 1.620 2.060 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.560 2.350 3.150 2.650 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.760 2.460 2.160 3.180 ;
        RECT  2.160 2.940 2.180 3.180 ;
        RECT  2.180 2.940 2.420 3.210 ;
        RECT  2.420 2.950 2.440 3.210 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.190 5.440 ;
        RECT  0.190 4.480 0.590 5.440 ;
        RECT  0.590 4.640 2.750 5.440 ;
        RECT  2.750 4.480 3.150 5.440 ;
        RECT  3.150 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        RECT  0.990 -0.400 1.390 0.560 ;
        RECT  1.390 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.570 1.220 3.730 1.460 ;
        RECT  3.330 0.800 3.570 1.460 ;
        RECT  2.210 0.800 3.330 1.040 ;
        RECT  1.970 0.800 2.210 1.540 ;
        RECT  1.810 1.140 1.970 1.540 ;
        RECT  0.570 1.220 1.810 1.460 ;
        RECT  0.170 1.140 0.570 1.540 ;
    END
END OAI22X1

MACRO OAI222XL
    CLASS CORE ;
    FOREIGN OAI222XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.770 3.540 2.190 3.940 ;
        RECT  4.450 1.270 4.610 1.670 ;
        RECT  2.190 3.700 4.700 3.940 ;
        RECT  4.610 1.270 4.850 2.100 ;
        RECT  4.700 3.700 5.100 4.100 ;
        RECT  5.100 3.700 5.170 4.060 ;
        RECT  5.170 3.700 5.480 4.020 ;
        RECT  5.480 3.510 5.490 4.020 ;
        RECT  4.850 1.860 5.490 2.100 ;
        RECT  5.490 1.860 5.730 4.020 ;
        RECT  5.730 3.510 5.740 3.770 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.410 2.940 4.170 3.360 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 2.380 4.720 2.660 ;
        RECT  4.720 2.380 4.950 2.790 ;
        RECT  4.950 2.390 5.120 2.790 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.220 2.650 ;
        RECT  0.220 2.390 0.460 3.110 ;
        RECT  0.460 2.660 0.550 3.110 ;
        RECT  0.550 2.710 0.920 3.110 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.820 1.250 2.100 ;
        RECT  1.250 1.820 1.650 2.320 ;
        RECT  1.650 1.820 1.660 2.100 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.390 3.100 2.650 ;
        RECT  3.100 2.390 3.170 2.630 ;
        RECT  3.170 2.210 3.570 2.630 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.940 2.010 3.220 ;
        RECT  2.010 2.700 2.410 3.220 ;
        RECT  2.410 2.940 2.420 3.220 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.480 5.440 ;
        RECT  0.480 4.480 0.880 5.440 ;
        RECT  0.880 4.640 3.220 5.440 ;
        RECT  3.220 4.480 3.620 5.440 ;
        RECT  3.620 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 1.780 0.560 ;
        RECT  1.780 -0.400 5.940 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.460 1.180 5.620 1.580 ;
        RECT  5.220 0.700 5.460 1.580 ;
        RECT  4.090 0.700 5.220 0.940 ;
        RECT  3.690 0.700 4.090 1.580 ;
        RECT  2.510 0.700 3.690 0.940 ;
        RECT  2.930 1.230 3.330 1.630 ;
        RECT  0.770 1.300 2.930 1.540 ;
        RECT  2.190 0.700 2.510 0.950 ;
        RECT  2.110 0.710 2.190 0.950 ;
    END
END OAI222XL

MACRO OAI222X4
    CLASS CORE ;
    FOREIGN OAI222X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI222XL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  7.250 1.100 7.260 1.500 ;
        RECT  7.260 1.090 7.360 1.500 ;
        RECT  7.250 3.180 7.370 3.580 ;
        RECT  7.360 1.090 7.370 2.710 ;
        RECT  7.370 1.090 7.390 3.580 ;
        RECT  7.390 1.090 7.740 3.590 ;
        RECT  7.740 1.820 7.810 3.590 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 2.950 3.650 3.210 ;
        RECT  3.650 2.750 3.760 3.210 ;
        RECT  3.760 2.750 4.050 3.200 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.610 2.290 5.010 2.690 ;
        RECT  5.010 2.290 5.070 2.650 ;
        RECT  5.070 2.390 5.080 2.650 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.950 0.460 3.220 ;
        RECT  0.460 2.960 0.820 3.220 ;
        RECT  0.820 2.760 1.220 3.220 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.820 1.450 2.100 ;
        RECT  1.450 1.820 1.850 2.330 ;
        RECT  1.850 1.820 1.860 2.100 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 1.830 3.190 2.090 ;
        RECT  3.190 1.830 3.620 2.230 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 2.950 2.280 3.210 ;
        RECT  2.280 2.400 2.440 3.210 ;
        RECT  2.440 2.400 2.520 3.200 ;
        RECT  2.520 2.400 2.850 2.640 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.830 5.440 ;
        RECT  0.830 3.780 0.840 5.440 ;
        RECT  0.840 3.580 1.240 5.440 ;
        RECT  1.240 3.780 1.250 5.440 ;
        RECT  1.250 4.640 3.340 5.440 ;
        RECT  3.340 4.480 3.740 5.440 ;
        RECT  3.740 4.640 6.480 5.440 ;
        RECT  6.480 3.720 6.490 5.440 ;
        RECT  6.490 3.520 6.890 5.440 ;
        RECT  6.890 3.720 6.900 5.440 ;
        RECT  6.900 4.640 8.090 5.440 ;
        RECT  8.090 3.220 8.330 5.440 ;
        RECT  8.330 4.640 8.580 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 1.420 ;
        RECT  0.170 -0.400 0.570 1.540 ;
        RECT  0.570 -0.400 0.580 1.420 ;
        RECT  0.580 -0.400 1.640 0.400 ;
        RECT  1.640 -0.400 2.040 0.560 ;
        RECT  2.040 -0.400 6.480 0.400 ;
        RECT  6.480 -0.400 6.490 0.770 ;
        RECT  6.490 -0.400 6.890 0.970 ;
        RECT  6.890 -0.400 6.900 0.770 ;
        RECT  6.900 -0.400 8.000 0.400 ;
        RECT  8.000 -0.400 8.010 1.060 ;
        RECT  8.010 -0.400 8.410 1.260 ;
        RECT  8.410 -0.400 8.420 1.060 ;
        RECT  8.420 -0.400 8.580 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.930 1.990 7.090 2.390 ;
        RECT  6.690 1.240 6.930 3.140 ;
        RECT  6.130 1.240 6.690 1.480 ;
        RECT  6.200 2.900 6.690 3.140 ;
        RECT  5.680 1.770 6.370 2.170 ;
        RECT  5.960 2.900 6.200 3.890 ;
        RECT  5.730 0.840 6.130 1.480 ;
        RECT  5.730 3.490 5.960 3.890 ;
        RECT  5.440 1.770 5.680 3.210 ;
        RECT  4.790 1.770 5.440 2.010 ;
        RECT  5.030 2.970 5.440 3.210 ;
        RECT  4.790 2.970 5.030 3.890 ;
        RECT  4.550 1.220 4.790 2.010 ;
        RECT  4.630 3.490 4.790 3.890 ;
        RECT  2.460 3.650 4.630 3.890 ;
        RECT  4.390 1.220 4.550 1.620 ;
        RECT  0.930 1.300 3.370 1.540 ;
        RECT  2.060 3.490 2.460 3.890 ;
    END
END OAI222X4

MACRO OAI222X2
    CLASS CORE ;
    FOREIGN OAI222X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI222XL ;
    SIZE 9.900 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.670 3.590 2.300 3.990 ;
        RECT  2.300 3.590 4.790 3.830 ;
        RECT  4.790 3.590 5.190 3.990 ;
        RECT  7.180 1.420 7.340 1.820 ;
        RECT  7.340 1.420 7.580 2.110 ;
        RECT  5.190 3.590 7.620 3.830 ;
        RECT  7.620 3.590 8.020 3.990 ;
        RECT  7.580 1.870 8.620 2.110 ;
        RECT  8.620 1.260 9.020 2.110 ;
        RECT  8.020 3.590 9.450 3.830 ;
        RECT  9.440 2.390 9.450 2.650 ;
        RECT  9.020 1.870 9.450 2.110 ;
        RECT  9.450 1.870 9.690 3.830 ;
        RECT  9.690 2.390 9.700 2.650 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.690 2.390 6.900 2.970 ;
        RECT  6.900 2.390 7.140 3.310 ;
        RECT  7.140 3.070 8.830 3.310 ;
        RECT  8.830 2.560 9.070 3.310 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.430 2.390 7.730 2.790 ;
        RECT  7.730 2.380 8.330 2.790 ;
        RECT  8.330 2.380 8.400 2.680 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.690 2.530 1.090 3.210 ;
        RECT  1.090 2.950 1.120 3.210 ;
        RECT  1.120 2.950 2.530 3.190 ;
        RECT  2.530 2.940 2.630 3.190 ;
        RECT  2.630 2.540 2.870 3.190 ;
        RECT  2.870 2.540 3.030 2.940 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.450 1.950 1.520 2.500 ;
        RECT  1.520 1.830 1.780 2.500 ;
        RECT  1.780 2.100 1.850 2.500 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 2.940 3.810 3.220 ;
        RECT  3.810 2.540 3.970 3.220 ;
        RECT  3.970 2.540 4.210 3.310 ;
        RECT  4.210 3.070 5.980 3.310 ;
        RECT  5.980 2.560 6.220 3.310 ;
        RECT  6.220 2.560 6.380 2.960 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.730 2.380 5.220 2.800 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.380 5.440 ;
        RECT  0.380 3.930 0.390 5.440 ;
        RECT  0.390 3.730 0.790 5.440 ;
        RECT  0.790 3.930 0.800 5.440 ;
        RECT  0.800 4.640 2.950 5.440 ;
        RECT  2.950 4.480 3.350 5.440 ;
        RECT  3.350 4.640 6.110 5.440 ;
        RECT  6.110 4.480 6.510 5.440 ;
        RECT  6.510 4.640 8.920 5.440 ;
        RECT  8.920 4.480 9.320 5.440 ;
        RECT  9.320 4.640 9.900 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 1.090 ;
        RECT  0.170 -0.400 0.570 1.290 ;
        RECT  0.570 -0.400 0.580 1.090 ;
        RECT  0.580 -0.400 1.710 0.400 ;
        RECT  1.710 -0.400 2.830 0.560 ;
        RECT  2.830 -0.400 9.900 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  9.340 0.740 9.740 1.380 ;
        RECT  8.300 0.740 9.340 0.980 ;
        RECT  8.060 0.740 8.300 1.590 ;
        RECT  7.900 1.190 8.060 1.590 ;
        RECT  5.740 1.450 6.140 1.850 ;
        RECT  4.640 1.450 5.740 1.690 ;
        RECT  4.240 1.450 4.640 2.060 ;
        RECT  2.720 1.450 4.240 1.690 ;
        RECT  2.320 1.290 2.720 1.690 ;
        RECT  1.320 1.290 2.320 1.530 ;
        RECT  0.920 1.130 1.320 1.530 ;
    END
END OAI222X2

MACRO OAI222X1
    CLASS CORE ;
    FOREIGN OAI222X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI222XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.140 3.490 2.540 3.890 ;
        RECT  2.540 3.490 2.970 3.780 ;
        RECT  2.970 3.490 4.800 3.730 ;
        RECT  4.550 1.200 4.870 1.440 ;
        RECT  4.870 1.200 5.110 1.620 ;
        RECT  4.800 3.490 5.200 3.890 ;
        RECT  5.110 1.380 5.390 1.620 ;
        RECT  5.200 3.490 5.490 3.780 ;
        RECT  5.390 1.380 5.490 1.820 ;
        RECT  5.490 1.380 5.730 3.780 ;
        RECT  5.730 3.510 5.740 3.780 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.070 1.770 4.550 2.170 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.710 2.470 5.130 3.220 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.380 0.690 2.680 ;
        RECT  0.690 2.270 0.990 2.680 ;
        RECT  0.990 2.270 1.090 2.670 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 1.120 3.210 ;
        RECT  1.120 2.950 1.530 3.190 ;
        RECT  1.530 1.980 1.770 3.190 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.940 3.320 3.220 ;
        RECT  3.320 2.450 3.560 3.220 ;
        RECT  3.560 2.450 3.720 2.960 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 2.390 2.380 2.650 ;
        RECT  2.380 2.200 2.780 2.650 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.910 5.440 ;
        RECT  0.910 3.720 0.920 5.440 ;
        RECT  0.920 3.520 1.320 5.440 ;
        RECT  1.320 3.720 1.330 5.440 ;
        RECT  1.330 4.640 3.460 5.440 ;
        RECT  3.460 4.480 3.860 5.440 ;
        RECT  3.860 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 1.350 ;
        RECT  0.170 -0.400 0.570 1.550 ;
        RECT  0.570 -0.400 0.580 1.350 ;
        RECT  0.580 -0.400 1.680 0.400 ;
        RECT  1.680 -0.400 1.690 1.060 ;
        RECT  1.690 -0.400 2.090 1.180 ;
        RECT  2.090 -0.400 2.100 1.060 ;
        RECT  2.100 -0.400 5.940 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.440 0.670 5.680 1.100 ;
        RECT  4.190 0.670 5.440 0.910 ;
        RECT  3.950 0.670 4.190 1.450 ;
        RECT  3.790 1.210 3.950 1.450 ;
        RECT  3.030 1.350 3.430 1.750 ;
        RECT  1.330 1.460 3.030 1.700 ;
        RECT  0.930 1.200 1.330 1.700 ;
    END
END OAI222X1

MACRO OAI221XL
    CLASS CORE ;
    FOREIGN OAI221XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.690 3.510 2.190 3.920 ;
        RECT  2.190 3.510 3.750 3.750 ;
        RECT  3.750 3.510 3.790 3.760 ;
        RECT  4.160 1.270 4.170 1.530 ;
        RECT  3.790 3.510 4.190 3.910 ;
        RECT  4.170 1.270 4.420 1.680 ;
        RECT  4.190 3.510 4.510 3.750 ;
        RECT  4.510 3.500 4.670 3.750 ;
        RECT  4.420 1.280 4.670 1.680 ;
        RECT  4.670 1.280 4.910 3.750 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 2.940 3.990 3.240 ;
        RECT  3.990 2.830 4.390 3.230 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.210 2.650 ;
        RECT  0.210 2.060 0.460 2.650 ;
        RECT  0.460 2.060 0.870 2.470 ;
        RECT  0.870 2.070 1.110 2.470 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.940 1.430 3.220 ;
        RECT  1.430 2.630 1.830 3.220 ;
        RECT  1.830 2.940 1.840 3.220 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.380 3.330 2.660 ;
        RECT  3.330 2.110 3.580 2.660 ;
        RECT  3.580 2.110 3.730 2.510 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.820 2.240 2.100 ;
        RECT  2.240 1.820 2.480 2.350 ;
        RECT  2.480 1.820 2.490 2.100 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.460 5.440 ;
        RECT  0.460 3.690 0.470 5.440 ;
        RECT  0.470 3.490 0.870 5.440 ;
        RECT  0.870 3.690 0.880 5.440 ;
        RECT  0.880 4.640 2.970 5.440 ;
        RECT  2.970 4.480 3.370 5.440 ;
        RECT  3.370 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 1.320 ;
        RECT  0.170 -0.400 0.570 1.520 ;
        RECT  0.570 -0.400 0.580 1.320 ;
        RECT  0.580 -0.400 1.740 0.400 ;
        RECT  1.740 -0.400 2.140 0.560 ;
        RECT  2.140 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.090 1.260 3.490 1.660 ;
        RECT  1.330 1.260 3.090 1.500 ;
        RECT  0.930 1.150 1.330 1.550 ;
    END
END OAI221XL

MACRO OAI221X4
    CLASS CORE ;
    FOREIGN OAI221X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI221XL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.580 2.800 6.590 3.770 ;
        RECT  6.590 2.800 6.710 4.260 ;
        RECT  6.590 1.270 6.710 1.670 ;
        RECT  6.710 1.260 6.990 4.260 ;
        RECT  6.990 1.260 7.000 3.770 ;
        RECT  7.000 1.260 7.130 3.220 ;
        RECT  7.130 1.820 7.150 3.220 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.820 3.850 2.100 ;
        RECT  3.850 1.820 4.090 2.530 ;
        RECT  4.090 2.130 4.250 2.530 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.360 2.650 ;
        RECT  0.360 2.060 0.460 2.650 ;
        RECT  0.460 2.060 0.600 2.630 ;
        RECT  0.600 2.060 0.670 2.470 ;
        RECT  0.670 2.070 0.920 2.470 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.940 1.290 3.220 ;
        RECT  1.290 2.710 1.690 3.220 ;
        RECT  1.690 2.940 1.700 3.220 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.950 2.950 3.210 ;
        RECT  2.950 2.620 3.100 3.210 ;
        RECT  3.100 2.620 3.120 3.190 ;
        RECT  3.120 2.460 3.190 3.190 ;
        RECT  3.190 2.460 3.520 2.860 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.120 2.090 2.600 2.660 ;
        RECT  2.600 2.100 2.660 2.660 ;
        RECT  2.660 2.320 2.670 2.660 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.320 5.440 ;
        RECT  0.320 3.750 0.330 5.440 ;
        RECT  0.330 3.550 0.730 5.440 ;
        RECT  0.730 3.750 0.740 5.440 ;
        RECT  0.740 4.640 2.830 5.440 ;
        RECT  2.830 4.480 3.230 5.440 ;
        RECT  3.230 4.640 5.820 5.440 ;
        RECT  5.820 3.870 5.830 5.440 ;
        RECT  5.830 3.670 6.230 5.440 ;
        RECT  6.230 3.870 6.240 5.440 ;
        RECT  6.240 4.640 7.340 5.440 ;
        RECT  7.340 4.080 7.350 5.440 ;
        RECT  7.350 3.880 7.750 5.440 ;
        RECT  7.750 4.080 7.760 5.440 ;
        RECT  7.760 4.640 7.920 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.380 0.400 ;
        RECT  1.380 -0.400 1.780 0.560 ;
        RECT  1.780 -0.400 5.820 0.400 ;
        RECT  5.820 -0.400 5.830 1.120 ;
        RECT  5.830 -0.400 6.230 1.320 ;
        RECT  6.230 -0.400 6.240 1.120 ;
        RECT  6.240 -0.400 7.340 0.400 ;
        RECT  7.340 -0.400 7.350 0.790 ;
        RECT  7.350 -0.400 7.750 0.990 ;
        RECT  7.750 -0.400 7.760 0.790 ;
        RECT  7.760 -0.400 7.920 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.260 1.950 6.440 2.350 ;
        RECT  6.020 1.950 6.260 3.390 ;
        RECT  5.550 1.950 6.020 2.190 ;
        RECT  5.470 3.150 6.020 3.390 ;
        RECT  4.770 2.470 5.710 2.870 ;
        RECT  5.310 0.670 5.550 2.190 ;
        RECT  5.070 3.140 5.470 4.120 ;
        RECT  5.070 0.670 5.310 0.910 ;
        RECT  4.770 1.330 4.850 1.730 ;
        RECT  4.530 1.330 4.770 3.760 ;
        RECT  4.450 1.330 4.530 1.730 ;
        RECT  4.060 3.520 4.530 3.760 ;
        RECT  3.860 3.520 4.060 3.920 ;
        RECT  3.870 1.040 4.030 1.440 ;
        RECT  3.630 0.680 3.870 1.440 ;
        RECT  1.750 3.510 3.860 3.930 ;
        RECT  2.510 0.680 3.630 0.920 ;
        RECT  3.110 1.210 3.270 1.450 ;
        RECT  2.870 1.210 3.110 1.820 ;
        RECT  1.830 1.580 2.870 1.820 ;
        RECT  2.270 0.680 2.510 1.300 ;
        RECT  2.110 1.060 2.270 1.300 ;
        RECT  1.590 1.270 1.830 1.820 ;
        RECT  1.550 3.520 1.750 3.920 ;
        RECT  1.170 1.270 1.590 1.510 ;
        RECT  0.770 1.110 1.170 1.510 ;
    END
END OAI221X4

MACRO OAI221X2
    CLASS CORE ;
    FOREIGN OAI221X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI221XL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.390 3.570 1.790 3.970 ;
        RECT  1.790 3.650 3.830 3.890 ;
        RECT  3.830 3.650 4.230 4.050 ;
        RECT  4.230 3.650 5.480 3.890 ;
        RECT  5.480 3.510 5.490 3.890 ;
        RECT  5.490 3.490 6.040 3.890 ;
        RECT  6.040 3.000 6.280 3.890 ;
        RECT  5.980 1.460 6.380 1.920 ;
        RECT  6.280 3.000 6.760 3.240 ;
        RECT  6.380 1.680 6.760 1.920 ;
        RECT  6.760 1.680 7.000 3.240 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.000 2.320 6.490 2.720 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.400 2.860 0.800 3.260 ;
        RECT  0.800 2.950 1.120 3.260 ;
        RECT  1.120 3.020 2.230 3.260 ;
        RECT  2.230 2.400 2.470 3.260 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 2.250 1.870 2.660 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.870 2.850 3.270 3.250 ;
        RECT  3.270 2.850 3.350 3.170 ;
        RECT  3.350 2.390 3.590 3.170 ;
        RECT  3.590 2.390 3.760 2.650 ;
        RECT  3.760 2.390 4.900 2.630 ;
        RECT  4.900 2.390 5.140 3.060 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.880 2.920 4.570 3.360 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.140 0.170 5.440 ;
        RECT  0.170 3.940 0.570 5.440 ;
        RECT  0.570 4.140 0.580 5.440 ;
        RECT  0.580 4.640 2.600 5.440 ;
        RECT  2.600 4.370 2.610 5.440 ;
        RECT  2.610 4.170 3.010 5.440 ;
        RECT  3.010 4.370 3.020 5.440 ;
        RECT  3.020 4.640 5.050 5.440 ;
        RECT  5.050 4.370 5.060 5.440 ;
        RECT  5.060 4.170 5.460 5.440 ;
        RECT  5.460 4.370 5.470 5.440 ;
        RECT  5.470 4.640 6.630 5.440 ;
        RECT  6.630 3.870 6.640 5.440 ;
        RECT  6.640 3.670 7.040 5.440 ;
        RECT  7.040 3.870 7.050 5.440 ;
        RECT  7.050 4.640 7.260 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 1.230 ;
        RECT  0.170 -0.400 0.570 1.430 ;
        RECT  0.570 -0.400 0.580 1.230 ;
        RECT  0.580 -0.400 1.680 0.400 ;
        RECT  1.680 -0.400 1.690 1.090 ;
        RECT  1.690 -0.400 2.090 1.290 ;
        RECT  2.090 -0.400 2.100 1.090 ;
        RECT  2.100 -0.400 3.200 0.400 ;
        RECT  3.200 -0.400 3.210 1.090 ;
        RECT  3.210 -0.400 3.610 1.290 ;
        RECT  3.610 -0.400 3.620 1.090 ;
        RECT  3.620 -0.400 7.260 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  7.090 0.920 7.100 1.320 ;
        RECT  6.700 0.900 7.090 1.320 ;
        RECT  5.590 0.900 6.700 1.140 ;
        RECT  5.190 0.670 5.590 1.140 ;
        RECT  3.950 0.670 5.190 0.910 ;
        RECT  4.560 1.580 4.960 2.060 ;
        RECT  2.850 1.580 4.560 1.820 ;
        RECT  2.450 1.350 2.850 1.820 ;
        RECT  1.330 1.580 2.450 1.820 ;
        RECT  0.930 1.350 1.330 1.820 ;
    END
END OAI221X2

MACRO OAI221X1
    CLASS CORE ;
    FOREIGN OAI221X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI221XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 3.490 1.920 3.890 ;
        RECT  1.920 3.490 2.310 3.780 ;
        RECT  2.310 3.520 4.260 3.760 ;
        RECT  4.260 3.330 4.730 3.760 ;
        RECT  4.730 3.220 4.790 3.760 ;
        RECT  4.630 1.130 4.790 1.530 ;
        RECT  4.790 1.130 4.820 3.760 ;
        RECT  4.820 1.130 5.030 3.770 ;
        RECT  5.030 3.510 5.080 3.770 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.000 2.550 4.080 2.950 ;
        RECT  4.080 2.400 4.160 2.950 ;
        RECT  4.160 2.390 4.400 2.950 ;
        RECT  4.400 2.390 4.420 2.650 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.060 0.430 2.650 ;
        RECT  0.430 2.050 0.460 2.650 ;
        RECT  0.460 2.050 0.680 2.450 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 0.970 3.210 ;
        RECT  0.970 2.630 1.120 3.210 ;
        RECT  1.120 2.630 1.210 3.190 ;
        RECT  1.210 2.630 1.640 3.090 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.950 2.860 3.210 ;
        RECT  2.860 2.940 3.100 3.210 ;
        RECT  3.100 2.940 3.280 3.180 ;
        RECT  3.280 2.550 3.520 3.180 ;
        RECT  3.520 2.550 3.680 2.950 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.530 2.090 ;
        RECT  1.530 1.830 1.780 2.280 ;
        RECT  1.780 2.040 2.060 2.280 ;
        RECT  2.060 2.040 2.460 2.440 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.200 5.440 ;
        RECT  0.200 4.480 0.600 5.440 ;
        RECT  0.600 4.640 2.840 5.440 ;
        RECT  2.840 4.480 3.240 5.440 ;
        RECT  3.240 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 1.170 ;
        RECT  0.170 -0.400 0.570 1.370 ;
        RECT  0.570 -0.400 0.580 1.170 ;
        RECT  0.580 -0.400 1.810 0.400 ;
        RECT  1.810 -0.400 2.210 0.560 ;
        RECT  2.210 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.870 1.130 4.270 1.760 ;
        RECT  2.730 1.520 3.870 1.760 ;
        RECT  3.090 0.880 3.490 1.240 ;
        RECT  1.390 0.880 3.090 1.120 ;
        RECT  2.330 1.460 2.730 1.760 ;
        RECT  0.990 0.810 1.390 1.210 ;
    END
END OAI221X1

MACRO OAI21XL
    CLASS CORE ;
    FOREIGN OAI21XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.450 3.130 1.850 3.530 ;
        RECT  1.850 3.130 1.870 3.500 ;
        RECT  1.870 3.130 2.840 3.370 ;
        RECT  2.840 2.950 2.850 3.370 ;
        RECT  2.510 1.180 2.850 1.580 ;
        RECT  2.850 1.180 2.910 3.370 ;
        RECT  2.910 1.280 3.090 3.370 ;
        RECT  3.090 2.950 3.100 3.210 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.110 2.370 2.190 2.770 ;
        RECT  2.180 1.830 2.190 2.090 ;
        RECT  2.190 1.830 2.430 2.770 ;
        RECT  2.430 1.830 2.440 2.090 ;
        RECT  2.430 2.370 2.510 2.770 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.460 2.420 ;
        RECT  0.460 1.990 0.870 2.420 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.230 1.900 1.390 2.300 ;
        RECT  1.390 1.900 1.520 2.630 ;
        RECT  1.520 1.900 1.630 2.650 ;
        RECT  1.630 2.390 1.780 2.650 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 2.270 5.440 ;
        RECT  2.270 4.480 2.670 5.440 ;
        RECT  2.670 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        RECT  0.980 -0.400 1.380 0.560 ;
        RECT  1.380 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  0.170 1.310 2.150 1.550 ;
    END
END OAI21XL

MACRO OAI21X4
    CLASS CORE ;
    FOREIGN OAI21X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI21XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.630 3.440 2.300 3.850 ;
        RECT  2.300 3.440 4.070 3.840 ;
        RECT  4.070 2.940 4.470 3.840 ;
        RECT  4.470 2.940 4.730 3.780 ;
        RECT  4.730 2.380 5.090 3.780 ;
        RECT  5.090 1.360 5.170 3.780 ;
        RECT  5.170 1.360 5.490 3.340 ;
        RECT  5.490 1.360 5.570 1.760 ;
        RECT  5.490 2.940 5.950 3.340 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.770 2.240 6.050 2.640 ;
        RECT  6.050 1.950 6.140 2.640 ;
        RECT  6.140 1.830 6.170 2.640 ;
        RECT  6.170 1.830 6.380 2.480 ;
        RECT  6.380 1.830 6.400 2.090 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.550 2.190 0.710 2.590 ;
        RECT  0.710 2.190 0.860 3.170 ;
        RECT  0.860 2.190 0.950 3.210 ;
        RECT  0.950 2.930 1.120 3.210 ;
        RECT  1.120 2.930 2.950 3.170 ;
        RECT  2.950 2.520 2.960 3.170 ;
        RECT  2.960 2.350 3.280 3.170 ;
        RECT  3.280 2.350 3.290 2.950 ;
        RECT  3.290 2.350 3.360 2.590 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 2.030 1.520 2.430 ;
        RECT  1.520 2.030 1.780 2.650 ;
        RECT  1.780 2.030 1.800 2.640 ;
        RECT  1.800 2.030 1.880 2.430 ;
        RECT  1.880 2.110 2.330 2.350 ;
        RECT  2.330 1.830 2.570 2.350 ;
        RECT  2.570 1.830 2.970 2.100 ;
        RECT  2.970 1.830 3.670 2.070 ;
        RECT  3.670 1.830 3.890 2.320 ;
        RECT  3.890 1.830 3.910 2.660 ;
        RECT  3.910 2.080 4.290 2.660 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.400 5.440 ;
        RECT  0.400 3.690 0.410 5.440 ;
        RECT  0.410 3.490 0.810 5.440 ;
        RECT  0.810 3.690 0.820 5.440 ;
        RECT  0.820 4.640 2.840 5.440 ;
        RECT  2.840 4.240 2.850 5.440 ;
        RECT  2.850 4.120 3.250 5.440 ;
        RECT  3.250 4.240 3.260 5.440 ;
        RECT  3.260 4.640 4.670 5.440 ;
        RECT  4.670 4.300 4.680 5.440 ;
        RECT  4.680 4.100 5.080 5.440 ;
        RECT  5.080 4.300 5.090 5.440 ;
        RECT  5.090 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.850 0.400 ;
        RECT  0.850 -0.400 0.860 1.040 ;
        RECT  0.860 -0.400 1.260 1.160 ;
        RECT  1.260 -0.400 1.270 1.040 ;
        RECT  1.270 -0.400 2.340 0.400 ;
        RECT  2.340 -0.400 2.740 0.560 ;
        RECT  2.740 -0.400 3.740 0.400 ;
        RECT  3.740 -0.400 4.140 0.560 ;
        RECT  4.140 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.810 0.720 6.240 0.960 ;
        RECT  4.570 0.720 4.810 1.630 ;
        RECT  4.410 1.230 4.570 1.630 ;
        RECT  1.970 1.310 4.410 1.550 ;
        RECT  1.650 1.310 1.970 1.700 ;
        RECT  0.570 1.460 1.650 1.700 ;
        RECT  0.170 1.380 0.570 1.780 ;
    END
END OAI21X4

MACRO OAI21X2
    CLASS CORE ;
    FOREIGN OAI21X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI21XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.420 3.580 1.000 3.980 ;
        RECT  1.000 3.580 2.980 3.820 ;
        RECT  2.980 3.580 3.380 3.980 ;
        RECT  3.910 1.230 4.070 1.630 ;
        RECT  3.380 3.580 4.170 3.820 ;
        RECT  4.160 2.950 4.170 3.210 ;
        RECT  4.170 2.950 4.180 3.820 ;
        RECT  4.070 1.230 4.180 1.980 ;
        RECT  4.180 1.230 4.310 3.820 ;
        RECT  4.310 1.740 4.420 3.820 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.410 2.260 3.900 2.660 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 2.250 2.410 2.650 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.660 2.500 1.060 3.210 ;
        RECT  1.060 2.950 1.120 3.210 ;
        RECT  1.120 2.950 2.530 3.190 ;
        RECT  2.530 2.940 2.740 3.190 ;
        RECT  2.740 2.260 2.980 3.190 ;
        RECT  2.980 2.260 3.140 2.660 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.700 5.440 ;
        RECT  1.700 4.480 2.100 5.440 ;
        RECT  2.100 4.640 3.800 5.440 ;
        RECT  3.800 4.480 4.200 5.440 ;
        RECT  4.200 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        RECT  0.980 -0.400 1.380 0.560 ;
        RECT  1.380 -0.400 2.380 0.400 ;
        RECT  2.380 -0.400 2.390 1.250 ;
        RECT  2.390 -0.400 2.790 1.450 ;
        RECT  2.790 -0.400 2.800 1.250 ;
        RECT  2.800 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.910 1.060 5.070 1.460 ;
        RECT  4.670 0.710 4.910 1.460 ;
        RECT  3.550 0.710 4.670 0.950 ;
        RECT  3.390 0.710 3.550 1.610 ;
        RECT  3.310 0.710 3.390 1.970 ;
        RECT  3.150 1.210 3.310 1.970 ;
        RECT  2.030 1.730 3.150 1.970 ;
        RECT  1.790 1.220 2.030 1.970 ;
        RECT  1.630 1.220 1.790 1.620 ;
        RECT  0.570 1.300 1.630 1.540 ;
        RECT  0.170 1.220 0.570 1.620 ;
    END
END OAI21X2

MACRO OAI21X1
    CLASS CORE ;
    FOREIGN OAI21X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI21XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.810 2.960 2.210 3.540 ;
        RECT  2.210 2.960 2.840 3.200 ;
        RECT  2.840 2.950 2.850 3.210 ;
        RECT  2.570 1.060 2.850 1.460 ;
        RECT  2.850 1.060 3.090 3.210 ;
        RECT  3.090 2.950 3.100 3.210 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.050 2.080 2.180 2.480 ;
        RECT  2.180 2.080 2.440 2.650 ;
        RECT  2.440 2.080 2.450 2.480 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.060 0.820 2.650 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.940 1.280 3.220 ;
        RECT  1.280 1.790 1.520 3.220 ;
        RECT  1.520 2.940 1.530 3.220 ;
        RECT  1.520 1.790 1.680 2.190 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.560 5.440 ;
        RECT  0.560 3.480 0.980 5.440 ;
        RECT  0.980 4.640 2.630 5.440 ;
        RECT  2.630 4.480 3.030 5.440 ;
        RECT  3.030 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        RECT  0.980 -0.400 0.990 0.680 ;
        RECT  0.990 -0.400 1.390 0.880 ;
        RECT  1.390 -0.400 1.400 0.680 ;
        RECT  1.400 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.810 1.060 2.210 1.460 ;
        RECT  0.570 1.160 1.810 1.400 ;
        RECT  0.170 1.060 0.570 1.460 ;
    END
END OAI21X1

MACRO OAI211XL
    CLASS CORE ;
    FOREIGN OAI211XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.650 2.960 2.050 3.360 ;
        RECT  2.050 2.960 2.190 3.280 ;
        RECT  2.190 3.040 2.970 3.280 ;
        RECT  3.060 1.030 3.270 1.430 ;
        RECT  2.970 2.950 3.390 3.280 ;
        RECT  3.390 2.950 3.500 3.760 ;
        RECT  3.500 2.950 3.550 3.770 ;
        RECT  3.270 1.020 3.550 1.430 ;
        RECT  3.550 1.020 3.760 3.770 ;
        RECT  3.760 1.020 3.790 3.760 ;
        RECT  3.790 1.020 3.800 1.520 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.090 2.200 2.510 2.680 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.750 1.700 3.270 2.100 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.060 0.500 2.670 ;
        RECT  0.500 2.060 0.800 2.470 ;
        RECT  0.800 2.070 0.850 2.470 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 1.120 3.210 ;
        RECT  1.120 2.950 1.130 3.190 ;
        RECT  1.130 2.230 1.370 3.190 ;
        RECT  1.370 2.230 1.390 2.470 ;
        RECT  1.390 2.070 1.790 2.470 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.370 5.440 ;
        RECT  0.370 4.480 0.770 5.440 ;
        RECT  0.770 4.640 2.480 5.440 ;
        RECT  2.480 4.480 2.880 5.440 ;
        RECT  2.880 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.000 0.400 ;
        RECT  1.000 -0.400 1.400 0.560 ;
        RECT  1.400 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.840 1.030 2.240 1.430 ;
        RECT  0.570 1.110 1.840 1.350 ;
        RECT  0.170 1.030 0.570 1.430 ;
    END
END OAI211XL

MACRO OAI211X4
    CLASS CORE ;
    FOREIGN OAI211X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI211XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.850 2.800 4.860 3.720 ;
        RECT  4.860 2.800 5.260 4.210 ;
        RECT  5.260 2.800 5.270 3.720 ;
        RECT  5.270 2.800 5.340 3.220 ;
        RECT  5.210 1.040 5.340 1.450 ;
        RECT  5.340 1.040 5.740 3.220 ;
        RECT  5.740 1.820 5.830 3.220 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.820 1.780 2.220 2.180 ;
        RECT  2.220 1.830 2.440 2.090 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.600 2.370 3.000 2.770 ;
        RECT  3.000 2.390 3.100 2.650 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 1.100 3.210 ;
        RECT  1.100 2.360 1.120 3.210 ;
        RECT  1.120 2.360 1.340 3.200 ;
        RECT  1.340 2.360 1.500 2.760 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.210 2.650 ;
        RECT  0.210 2.390 0.360 2.670 ;
        RECT  0.360 2.360 0.810 2.680 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.450 5.440 ;
        RECT  1.450 4.480 2.990 5.440 ;
        RECT  2.990 4.640 4.090 5.440 ;
        RECT  4.090 4.350 4.100 5.440 ;
        RECT  4.100 4.150 4.500 5.440 ;
        RECT  4.500 4.350 4.510 5.440 ;
        RECT  4.510 4.640 5.690 5.440 ;
        RECT  5.690 3.840 5.700 5.440 ;
        RECT  5.700 3.640 6.100 5.440 ;
        RECT  6.100 3.840 6.110 5.440 ;
        RECT  6.110 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.880 0.400 ;
        RECT  0.880 -0.400 1.280 0.560 ;
        RECT  1.280 -0.400 4.390 0.400 ;
        RECT  4.390 -0.400 4.790 0.560 ;
        RECT  4.790 -0.400 6.000 0.400 ;
        RECT  6.000 -0.400 6.010 0.850 ;
        RECT  6.010 -0.400 6.410 1.050 ;
        RECT  6.410 -0.400 6.420 0.850 ;
        RECT  6.420 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.580 2.120 5.020 2.520 ;
        RECT  4.340 1.130 4.580 3.860 ;
        RECT  3.970 1.130 4.340 1.370 ;
        RECT  3.740 3.620 4.340 3.860 ;
        RECT  3.700 2.030 4.060 2.430 ;
        RECT  3.570 0.970 3.970 1.370 ;
        RECT  3.340 3.620 3.740 4.020 ;
        RECT  3.460 1.650 3.700 3.340 ;
        RECT  3.210 1.650 3.460 1.890 ;
        RECT  2.600 3.100 3.460 3.340 ;
        RECT  2.970 1.100 3.210 1.890 ;
        RECT  2.810 1.100 2.970 1.500 ;
        RECT  2.440 3.100 2.600 3.600 ;
        RECT  2.200 3.100 2.440 3.940 ;
        RECT  0.580 3.700 2.200 3.940 ;
        RECT  1.590 1.100 1.990 1.500 ;
        RECT  0.570 1.160 1.590 1.400 ;
        RECT  0.180 3.700 0.580 4.130 ;
        RECT  0.170 1.050 0.570 1.450 ;
    END
END OAI211X4

MACRO OAI211X2
    CLASS CORE ;
    FOREIGN OAI211X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI211XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.530 3.610 0.930 4.010 ;
        RECT  0.930 3.610 3.090 3.850 ;
        RECT  3.090 3.610 3.490 4.030 ;
        RECT  3.490 3.610 4.610 3.850 ;
        RECT  4.550 1.360 4.950 1.850 ;
        RECT  4.610 3.610 5.010 4.030 ;
        RECT  5.010 3.610 6.150 3.850 ;
        RECT  6.140 2.390 6.150 2.650 ;
        RECT  4.950 1.610 6.150 1.850 ;
        RECT  6.150 1.610 6.390 3.850 ;
        RECT  6.390 2.390 6.400 2.650 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.720 2.940 3.730 3.220 ;
        RECT  3.570 2.230 3.730 2.630 ;
        RECT  3.730 2.230 3.970 3.220 ;
        RECT  3.970 2.940 5.350 3.220 ;
        RECT  5.350 2.930 5.750 3.330 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.370 2.240 4.770 2.650 ;
        RECT  4.770 2.390 5.080 2.650 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.500 2.070 1.520 2.470 ;
        RECT  1.520 2.070 1.780 2.650 ;
        RECT  1.780 2.070 2.480 2.470 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.760 2.470 0.860 3.200 ;
        RECT  0.860 2.470 1.120 3.210 ;
        RECT  1.120 2.470 1.160 3.170 ;
        RECT  1.160 2.930 2.810 3.170 ;
        RECT  2.810 2.310 2.850 3.170 ;
        RECT  2.850 2.230 3.050 3.170 ;
        RECT  3.050 2.230 3.250 2.630 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.810 5.440 ;
        RECT  1.810 4.480 2.210 5.440 ;
        RECT  2.210 4.640 3.840 5.440 ;
        RECT  3.840 4.330 3.850 5.440 ;
        RECT  3.850 4.130 4.250 5.440 ;
        RECT  4.250 4.330 4.260 5.440 ;
        RECT  4.260 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        RECT  0.990 -0.400 1.390 0.560 ;
        RECT  1.390 -0.400 2.560 0.400 ;
        RECT  2.560 -0.400 2.570 1.060 ;
        RECT  2.570 -0.400 2.970 1.260 ;
        RECT  2.970 -0.400 2.980 1.060 ;
        RECT  2.980 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.770 0.840 6.170 1.320 ;
        RECT  3.730 0.840 5.770 1.080 ;
        RECT  3.570 0.840 3.730 1.520 ;
        RECT  3.490 0.840 3.570 1.790 ;
        RECT  3.330 1.120 3.490 1.790 ;
        RECT  2.210 1.550 3.330 1.790 ;
        RECT  1.970 1.110 2.210 1.790 ;
        RECT  1.810 1.110 1.970 1.550 ;
        RECT  0.570 1.310 1.810 1.550 ;
        RECT  0.170 1.150 0.570 1.550 ;
    END
END OAI211X2

MACRO OAI211X1
    CLASS CORE ;
    FOREIGN OAI211X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ OAI211XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.500 3.250 1.900 3.650 ;
        RECT  1.900 3.330 2.190 3.650 ;
        RECT  2.190 3.330 3.260 3.570 ;
        RECT  2.990 1.100 3.500 1.510 ;
        RECT  3.260 3.170 3.510 3.570 ;
        RECT  3.500 1.100 3.510 1.530 ;
        RECT  3.510 1.100 3.750 3.570 ;
        RECT  3.750 1.100 3.760 1.530 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.630 2.090 ;
        RECT  1.630 1.830 1.780 2.100 ;
        RECT  1.780 1.840 1.870 2.100 ;
        RECT  1.870 1.860 2.020 2.100 ;
        RECT  2.020 1.860 2.260 2.570 ;
        RECT  2.260 2.170 2.420 2.570 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.740 1.840 2.840 2.330 ;
        RECT  2.840 1.830 3.100 2.330 ;
        RECT  3.100 1.930 3.140 2.330 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.550 2.420 ;
        RECT  0.550 2.010 0.920 2.410 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 0.970 3.210 ;
        RECT  0.970 2.690 1.120 3.210 ;
        RECT  1.120 2.690 1.210 3.190 ;
        RECT  1.210 2.690 1.260 2.930 ;
        RECT  1.260 2.370 1.500 2.930 ;
        RECT  1.500 2.370 1.660 2.770 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.270 5.440 ;
        RECT  0.270 3.690 0.280 5.440 ;
        RECT  0.280 3.490 0.680 5.440 ;
        RECT  0.680 3.690 0.690 5.440 ;
        RECT  0.690 4.640 2.320 5.440 ;
        RECT  2.320 4.480 2.720 5.440 ;
        RECT  2.720 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        RECT  0.980 -0.400 0.990 0.900 ;
        RECT  0.990 -0.400 1.390 1.020 ;
        RECT  1.390 -0.400 1.400 0.900 ;
        RECT  1.400 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.770 0.990 2.170 1.550 ;
        RECT  0.570 1.310 1.770 1.550 ;
        RECT  0.170 1.020 0.570 1.550 ;
    END
END OAI211X1

MACRO NOR4BBXL
    CLASS CORE ;
    FOREIGN NOR4BBXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.710 1.280 3.080 1.520 ;
        RECT  3.080 1.260 3.410 1.520 ;
        RECT  3.410 0.860 3.650 1.520 ;
        RECT  3.420 3.510 3.820 3.930 ;
        RECT  3.650 0.860 3.850 1.280 ;
        RECT  3.850 0.860 4.820 1.100 ;
        RECT  4.820 0.710 5.080 1.100 ;
        RECT  3.820 3.690 5.540 3.930 ;
        RECT  5.080 0.860 5.540 1.100 ;
        RECT  5.540 0.860 5.780 3.930 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.370 2.420 1.610 3.210 ;
        RECT  1.610 2.950 1.780 3.210 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.000 1.820 2.530 2.240 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 2.390 4.420 2.650 ;
        RECT  4.420 2.410 4.500 2.650 ;
        RECT  4.500 2.410 4.740 2.820 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.620 0.570 3.220 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.210 5.440 ;
        RECT  1.210 4.480 1.610 5.440 ;
        RECT  1.610 4.640 4.160 5.440 ;
        RECT  4.160 4.480 4.560 5.440 ;
        RECT  4.560 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 2.380 0.400 ;
        RECT  2.380 -0.400 2.780 0.560 ;
        RECT  2.780 -0.400 4.060 0.400 ;
        RECT  4.060 -0.400 4.460 0.560 ;
        RECT  4.460 -0.400 5.940 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.020 1.390 5.260 3.410 ;
        RECT  3.050 1.870 5.020 2.110 ;
        RECT  3.550 2.420 3.790 2.820 ;
        RECT  2.900 2.580 3.550 2.820 ;
        RECT  2.810 1.870 3.050 2.270 ;
        RECT  2.660 2.580 2.900 3.740 ;
        RECT  1.080 3.500 2.660 3.740 ;
        RECT  0.840 1.290 1.080 3.740 ;
        RECT  0.180 1.290 0.840 1.530 ;
        RECT  0.660 3.490 0.840 3.740 ;
        RECT  0.260 3.490 0.660 3.890 ;
    END
END NOR4BBXL

MACRO NOR4BBX4
    CLASS CORE ;
    FOREIGN NOR4BBX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR4BBXL ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.690 0.860 3.670 1.100 ;
        RECT  3.670 0.860 3.910 1.380 ;
        RECT  3.910 1.140 7.980 1.380 ;
        RECT  7.980 0.780 8.030 1.380 ;
        RECT  8.030 0.700 8.470 2.100 ;
        RECT  3.540 3.940 11.940 4.180 ;
        RECT  8.470 0.860 11.940 1.100 ;
        RECT  11.940 0.860 12.180 4.180 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.590 1.630 3.210 ;
        RECT  1.630 2.590 1.760 3.660 ;
        RECT  1.760 2.950 1.780 3.660 ;
        RECT  1.780 2.970 1.870 3.660 ;
        RECT  1.870 3.420 5.780 3.660 ;
        RECT  5.780 2.700 6.180 3.660 ;
        RECT  6.180 3.420 9.850 3.660 ;
        RECT  9.850 2.620 10.090 3.660 ;
        RECT  10.090 2.620 10.250 3.020 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.110 1.950 2.290 2.650 ;
        RECT  2.290 1.950 2.510 3.090 ;
        RECT  2.510 2.410 2.530 3.090 ;
        RECT  2.530 2.850 4.990 3.090 ;
        RECT  4.990 2.180 5.230 3.090 ;
        RECT  5.230 2.180 5.390 2.580 ;
        RECT  5.390 2.180 6.510 2.420 ;
        RECT  6.510 2.180 6.680 2.580 ;
        RECT  6.680 2.180 6.920 3.130 ;
        RECT  6.920 2.890 9.260 3.130 ;
        RECT  9.260 1.900 9.500 3.130 ;
        RECT  9.500 1.900 9.780 2.300 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  10.670 2.160 11.140 2.660 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.390 2.650 ;
        RECT  0.390 2.060 0.460 2.650 ;
        RECT  0.460 2.060 0.630 2.640 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.280 5.440 ;
        RECT  1.280 4.480 1.680 5.440 ;
        RECT  1.680 4.640 5.750 5.440 ;
        RECT  5.750 4.480 6.150 5.440 ;
        RECT  6.150 4.640 10.150 5.440 ;
        RECT  10.150 4.480 10.550 5.440 ;
        RECT  10.550 4.640 12.540 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.920 0.400 ;
        RECT  0.920 -0.400 0.930 0.820 ;
        RECT  0.930 -0.400 1.330 1.020 ;
        RECT  1.330 -0.400 1.340 0.820 ;
        RECT  1.340 -0.400 2.510 0.400 ;
        RECT  2.510 -0.400 2.910 0.560 ;
        RECT  2.910 -0.400 4.180 0.400 ;
        RECT  4.180 -0.400 4.190 0.740 ;
        RECT  4.190 -0.400 4.590 0.860 ;
        RECT  4.590 -0.400 4.600 0.740 ;
        RECT  4.600 -0.400 7.150 0.400 ;
        RECT  7.150 -0.400 7.160 0.740 ;
        RECT  7.160 -0.400 7.560 0.860 ;
        RECT  7.560 -0.400 7.570 0.740 ;
        RECT  7.570 -0.400 8.800 0.400 ;
        RECT  8.800 -0.400 9.040 0.560 ;
        RECT  9.040 -0.400 9.510 0.590 ;
        RECT  9.510 -0.400 10.440 0.400 ;
        RECT  10.440 -0.400 10.840 0.560 ;
        RECT  10.840 -0.400 12.540 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  11.420 1.380 11.660 3.490 ;
        RECT  8.980 1.380 11.420 1.620 ;
        RECT  11.370 3.250 11.420 3.490 ;
        RECT  10.970 3.250 11.370 3.650 ;
        RECT  8.740 1.380 8.980 2.610 ;
        RECT  7.630 2.370 8.740 2.610 ;
        RECT  7.470 2.170 7.630 2.610 ;
        RECT  7.230 1.660 7.470 2.610 ;
        RECT  4.670 1.660 7.230 1.900 ;
        RECT  4.430 1.660 4.670 2.570 ;
        RECT  4.270 2.170 4.430 2.570 ;
        RECT  3.230 2.330 4.270 2.570 ;
        RECT  3.940 1.810 3.950 2.050 ;
        RECT  3.550 1.730 3.940 2.050 ;
        RECT  3.140 1.730 3.550 1.970 ;
        RECT  2.830 2.250 3.230 2.570 ;
        RECT  2.900 1.380 3.140 1.970 ;
        RECT  1.160 1.380 2.900 1.620 ;
        RECT  0.920 1.310 1.160 3.780 ;
        RECT  0.570 1.310 0.920 1.550 ;
        RECT  0.770 3.540 0.920 3.780 ;
        RECT  0.370 3.540 0.770 3.940 ;
        RECT  0.170 1.060 0.570 1.550 ;
    END
END NOR4BBX4

MACRO NOR4BBX2
    CLASS CORE ;
    FOREIGN NOR4BBX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR4BBXL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.470 3.940 4.070 4.340 ;
        RECT  4.070 3.940 4.170 4.320 ;
        RECT  1.810 0.860 4.930 1.100 ;
        RECT  4.930 0.680 5.170 1.100 ;
        RECT  5.170 0.680 6.800 0.920 ;
        RECT  6.800 0.680 7.060 0.970 ;
        RECT  4.170 3.940 7.450 4.180 ;
        RECT  7.060 0.680 7.450 0.920 ;
        RECT  7.450 0.680 7.690 4.180 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.350 2.420 1.520 3.760 ;
        RECT  1.520 2.420 1.590 3.770 ;
        RECT  1.590 3.510 1.780 3.770 ;
        RECT  1.780 3.520 2.950 3.760 ;
        RECT  2.950 3.420 3.190 3.760 ;
        RECT  3.190 3.420 5.540 3.660 ;
        RECT  5.540 2.430 5.780 3.660 ;
        RECT  5.780 2.430 6.010 2.670 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.990 1.990 2.140 2.390 ;
        RECT  2.140 1.990 2.390 3.210 ;
        RECT  2.390 2.900 2.440 3.210 ;
        RECT  2.440 2.900 4.970 3.140 ;
        RECT  4.970 2.410 5.210 3.140 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.140 2.950 6.290 3.210 ;
        RECT  6.290 2.420 6.400 3.210 ;
        RECT  6.400 2.420 6.530 3.200 ;
        RECT  6.530 2.420 6.650 2.820 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.150 1.820 0.550 2.680 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.210 5.440 ;
        RECT  1.210 4.480 1.610 5.440 ;
        RECT  1.610 4.640 5.910 5.440 ;
        RECT  5.910 4.480 6.310 5.440 ;
        RECT  6.310 4.640 7.920 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.060 0.400 ;
        RECT  1.060 -0.400 1.480 1.020 ;
        RECT  1.480 -0.400 2.610 0.400 ;
        RECT  2.610 -0.400 3.010 0.560 ;
        RECT  3.010 -0.400 4.210 0.400 ;
        RECT  4.210 -0.400 4.610 0.560 ;
        RECT  4.610 -0.400 7.920 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.930 1.770 7.170 3.660 ;
        RECT  5.880 1.770 6.930 2.010 ;
        RECT  6.810 3.260 6.930 3.660 ;
        RECT  5.440 1.210 5.880 2.010 ;
        RECT  4.610 1.770 5.440 2.010 ;
        RECT  4.370 1.770 4.610 2.620 ;
        RECT  3.270 2.380 4.370 2.620 ;
        RECT  3.870 1.860 4.070 2.100 ;
        RECT  3.630 1.380 3.870 2.100 ;
        RECT  1.060 1.380 3.630 1.620 ;
        RECT  2.870 1.980 3.270 2.620 ;
        RECT  0.820 1.290 1.060 3.730 ;
        RECT  0.170 1.290 0.820 1.530 ;
        RECT  0.710 3.490 0.820 3.730 ;
        RECT  0.310 3.490 0.710 3.890 ;
    END
END NOR4BBX2

MACRO NOR4BBX1
    CLASS CORE ;
    FOREIGN NOR4BBX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR4BBXL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.740 1.230 3.390 1.470 ;
        RECT  3.390 0.860 3.630 1.470 ;
        RECT  3.420 3.510 3.820 3.950 ;
        RECT  3.630 0.860 4.820 1.100 ;
        RECT  4.820 0.710 5.080 1.100 ;
        RECT  3.820 3.710 5.540 3.950 ;
        RECT  5.080 0.860 5.540 1.100 ;
        RECT  5.540 0.860 5.780 3.950 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.370 2.420 1.610 3.210 ;
        RECT  1.610 2.950 1.780 3.210 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.000 1.830 2.400 2.260 ;
        RECT  2.400 1.830 2.440 2.090 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 2.390 4.420 2.650 ;
        RECT  4.420 2.410 4.500 2.650 ;
        RECT  4.500 2.410 4.740 2.820 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.570 2.420 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.210 5.440 ;
        RECT  1.210 4.480 1.610 5.440 ;
        RECT  1.610 4.640 4.160 5.440 ;
        RECT  4.160 4.480 4.560 5.440 ;
        RECT  4.560 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.130 0.400 ;
        RECT  1.130 -0.400 1.530 0.560 ;
        RECT  1.530 -0.400 2.420 0.400 ;
        RECT  2.420 -0.400 2.820 0.560 ;
        RECT  2.820 -0.400 4.050 0.400 ;
        RECT  4.050 -0.400 4.450 0.560 ;
        RECT  4.450 -0.400 5.940 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.020 1.390 5.260 3.430 ;
        RECT  3.040 1.870 5.020 2.110 ;
        RECT  3.560 2.420 3.800 2.820 ;
        RECT  2.900 2.580 3.560 2.820 ;
        RECT  2.800 1.870 3.040 2.270 ;
        RECT  2.660 2.580 2.900 3.730 ;
        RECT  1.080 3.490 2.660 3.730 ;
        RECT  0.840 1.310 1.080 3.730 ;
        RECT  0.260 1.310 0.840 1.550 ;
        RECT  0.670 3.490 0.840 3.730 ;
        RECT  0.270 3.490 0.670 3.890 ;
    END
END NOR4BBX1

MACRO NOR4BXL
    CLASS CORE ;
    FOREIGN NOR4BXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.410 3.530 3.810 3.930 ;
        RECT  3.810 3.530 4.170 3.770 ;
        RECT  4.160 2.950 4.170 3.210 ;
        RECT  1.820 1.290 4.170 1.530 ;
        RECT  4.170 1.290 4.410 3.770 ;
        RECT  4.410 2.950 4.420 3.210 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 2.660 1.930 3.210 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.990 1.800 2.450 2.200 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.820 2.140 3.190 2.650 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.570 2.420 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.210 5.440 ;
        RECT  1.210 4.480 1.610 5.440 ;
        RECT  1.610 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.130 0.400 ;
        RECT  1.130 -0.400 1.530 0.560 ;
        RECT  1.530 -0.400 2.520 0.400 ;
        RECT  2.520 -0.400 2.920 0.560 ;
        RECT  2.920 -0.400 4.060 0.400 ;
        RECT  4.060 -0.400 4.460 0.560 ;
        RECT  4.460 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.560 2.680 3.800 3.210 ;
        RECT  2.900 2.970 3.560 3.210 ;
        RECT  2.660 2.970 2.900 3.740 ;
        RECT  1.080 3.500 2.660 3.740 ;
        RECT  0.840 1.290 1.080 3.740 ;
        RECT  0.260 1.290 0.840 1.530 ;
        RECT  0.660 3.490 0.840 3.740 ;
        RECT  0.260 3.490 0.660 3.890 ;
    END
END NOR4BXL

MACRO NOR4BX4
    CLASS CORE ;
    FOREIGN NOR4BX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR4BXL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.690 0.750 1.740 1.150 ;
        RECT  1.740 0.750 2.090 1.160 ;
        RECT  2.090 0.860 3.320 1.160 ;
        RECT  3.430 3.890 3.480 4.290 ;
        RECT  3.480 3.880 3.830 4.290 ;
        RECT  3.320 0.860 3.990 1.390 ;
        RECT  3.990 0.970 4.820 1.390 ;
        RECT  3.830 3.880 8.070 4.180 ;
        RECT  8.070 3.880 8.910 4.340 ;
        RECT  4.820 0.960 9.680 1.390 ;
        RECT  9.680 0.960 10.360 1.550 ;
        RECT  8.910 3.880 10.670 4.180 ;
        RECT  10.360 0.970 10.670 1.550 ;
        RECT  10.670 0.970 10.970 4.180 ;
        RECT  10.970 0.970 11.090 3.220 ;
        RECT  11.090 1.820 11.110 3.220 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.950 1.530 3.210 ;
        RECT  1.530 2.590 1.630 3.210 ;
        RECT  1.630 2.590 1.770 3.610 ;
        RECT  1.770 2.950 1.780 3.610 ;
        RECT  1.780 2.970 1.870 3.610 ;
        RECT  1.870 3.370 5.780 3.610 ;
        RECT  5.780 2.700 6.180 3.610 ;
        RECT  6.180 3.370 9.990 3.610 ;
        RECT  9.990 2.620 10.230 3.610 ;
        RECT  10.230 2.620 10.390 3.020 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.930 1.950 2.090 2.190 ;
        RECT  2.090 1.950 2.180 2.630 ;
        RECT  2.180 1.950 2.290 2.650 ;
        RECT  2.290 1.950 2.330 3.050 ;
        RECT  2.330 2.390 2.440 3.050 ;
        RECT  2.440 2.410 2.530 3.050 ;
        RECT  2.530 2.810 4.980 3.050 ;
        RECT  4.980 2.180 5.220 3.050 ;
        RECT  5.220 2.180 5.380 2.580 ;
        RECT  5.380 2.180 6.510 2.420 ;
        RECT  6.510 2.180 6.680 2.580 ;
        RECT  6.680 2.180 6.920 3.010 ;
        RECT  6.920 2.770 9.450 3.010 ;
        RECT  9.450 1.900 9.690 3.010 ;
        RECT  9.690 1.900 9.910 2.300 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.800 2.250 3.200 2.570 ;
        RECT  3.200 2.330 4.270 2.570 ;
        RECT  4.270 2.170 4.430 2.570 ;
        RECT  4.430 1.660 4.670 2.570 ;
        RECT  4.670 1.660 7.300 1.900 ;
        RECT  7.300 1.660 7.540 2.490 ;
        RECT  7.540 1.650 7.810 2.490 ;
        RECT  7.810 2.250 9.070 2.490 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.390 2.650 ;
        RECT  0.390 2.060 0.460 2.650 ;
        RECT  0.460 2.060 0.630 2.640 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.170 5.440 ;
        RECT  1.170 4.480 1.570 5.440 ;
        RECT  1.570 4.640 5.750 5.440 ;
        RECT  5.750 4.480 6.150 5.440 ;
        RECT  6.150 4.640 10.270 5.440 ;
        RECT  10.270 4.480 10.670 5.440 ;
        RECT  10.670 4.640 11.880 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.920 0.400 ;
        RECT  0.920 -0.400 0.930 0.830 ;
        RECT  0.930 -0.400 1.330 1.030 ;
        RECT  1.330 -0.400 1.340 0.830 ;
        RECT  1.340 -0.400 2.510 0.400 ;
        RECT  2.510 -0.400 2.910 0.560 ;
        RECT  2.910 -0.400 4.150 0.400 ;
        RECT  4.150 -0.400 4.550 0.560 ;
        RECT  4.550 -0.400 7.330 0.400 ;
        RECT  7.330 -0.400 7.730 0.560 ;
        RECT  7.730 -0.400 8.970 0.400 ;
        RECT  8.970 -0.400 9.370 0.560 ;
        RECT  9.370 -0.400 10.610 0.400 ;
        RECT  10.610 -0.400 11.010 0.560 ;
        RECT  11.010 -0.400 11.880 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.540 1.660 3.940 2.050 ;
        RECT  2.950 1.660 3.540 1.900 ;
        RECT  2.710 1.430 2.950 1.900 ;
        RECT  1.160 1.430 2.710 1.670 ;
        RECT  0.920 1.310 1.160 3.780 ;
        RECT  0.570 1.310 0.920 1.550 ;
        RECT  0.740 3.540 0.920 3.780 ;
        RECT  0.340 3.540 0.740 3.940 ;
        RECT  0.170 1.060 0.570 1.550 ;
    END
END NOR4BX4

MACRO NOR4BX2
    CLASS CORE ;
    FOREIGN NOR4BX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR4BXL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.830 0.860 6.050 1.100 ;
        RECT  6.050 0.860 6.140 1.270 ;
        RECT  3.600 3.540 6.200 3.780 ;
        RECT  6.140 0.860 6.200 1.530 ;
        RECT  6.200 0.860 6.440 3.780 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.220 2.440 1.460 3.250 ;
        RECT  1.460 3.010 2.100 3.250 ;
        RECT  2.100 3.010 2.180 3.760 ;
        RECT  2.180 3.010 2.530 3.770 ;
        RECT  2.530 3.010 5.680 3.250 ;
        RECT  5.680 2.410 5.920 3.250 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.260 1.450 2.500 2.180 ;
        RECT  2.500 1.450 5.280 1.690 ;
        RECT  5.280 1.450 5.480 2.080 ;
        RECT  5.480 1.450 5.520 2.090 ;
        RECT  5.520 1.830 5.740 2.090 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.950 1.970 4.710 2.210 ;
        RECT  4.710 1.970 4.820 2.640 ;
        RECT  4.820 1.970 4.950 2.650 ;
        RECT  4.950 2.390 5.080 2.650 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 1.200 1.230 1.630 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.390 5.440 ;
        RECT  1.390 4.020 1.400 5.440 ;
        RECT  1.400 3.820 1.800 5.440 ;
        RECT  1.800 4.020 1.810 5.440 ;
        RECT  1.810 4.640 5.950 5.440 ;
        RECT  5.950 4.480 6.350 5.440 ;
        RECT  6.350 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.000 0.400 ;
        RECT  1.000 -0.400 1.010 0.410 ;
        RECT  1.010 -0.400 1.410 0.560 ;
        RECT  1.410 -0.400 1.420 0.410 ;
        RECT  1.420 -0.400 2.650 0.400 ;
        RECT  2.650 -0.400 3.050 0.560 ;
        RECT  3.050 -0.400 4.290 0.400 ;
        RECT  4.290 -0.400 4.690 0.560 ;
        RECT  4.690 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.970 2.490 4.110 2.730 ;
        RECT  1.730 1.900 1.970 2.730 ;
        RECT  0.400 1.900 1.730 2.140 ;
        RECT  0.400 0.670 0.570 0.910 ;
        RECT  0.400 3.010 0.570 3.990 ;
        RECT  0.170 0.670 0.400 3.990 ;
        RECT  0.160 0.670 0.170 3.980 ;
    END
END NOR4BX2

MACRO NOR4BX1
    CLASS CORE ;
    FOREIGN NOR4BX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR4BXL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.740 1.150 2.140 1.550 ;
        RECT  2.140 1.280 2.190 1.550 ;
        RECT  2.190 1.310 3.090 1.550 ;
        RECT  3.090 1.260 3.230 1.550 ;
        RECT  3.230 1.150 3.630 1.550 ;
        RECT  3.410 3.510 3.810 3.910 ;
        RECT  3.810 3.510 4.170 3.780 ;
        RECT  4.160 2.950 4.170 3.210 ;
        RECT  3.630 1.310 4.170 1.550 ;
        RECT  4.170 1.310 4.400 3.780 ;
        RECT  4.400 1.310 4.410 3.760 ;
        RECT  4.410 2.950 4.420 3.210 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.370 2.420 1.610 3.210 ;
        RECT  1.610 2.950 1.780 3.210 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.000 1.830 2.400 2.260 ;
        RECT  2.400 1.830 2.440 2.090 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.800 1.870 3.090 2.650 ;
        RECT  3.090 2.390 3.100 2.650 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.570 2.420 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.210 5.440 ;
        RECT  1.210 4.480 1.610 5.440 ;
        RECT  1.610 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.130 0.400 ;
        RECT  1.130 -0.400 1.530 0.560 ;
        RECT  1.530 -0.400 2.420 0.400 ;
        RECT  2.420 -0.400 2.820 0.560 ;
        RECT  2.820 -0.400 4.050 0.400 ;
        RECT  4.050 -0.400 4.450 0.560 ;
        RECT  4.450 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.560 2.430 3.800 3.210 ;
        RECT  2.900 2.970 3.560 3.210 ;
        RECT  2.660 2.970 2.900 3.740 ;
        RECT  1.080 3.500 2.660 3.740 ;
        RECT  0.840 1.320 1.080 3.740 ;
        RECT  0.260 1.320 0.840 1.560 ;
        RECT  0.670 3.500 0.840 3.740 ;
        RECT  0.270 3.500 0.670 3.960 ;
    END
END NOR4BX1

MACRO NOR4XL
    CLASS CORE ;
    FOREIGN NOR4XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.760 3.240 3.410 3.640 ;
        RECT  3.410 3.220 3.500 3.640 ;
        RECT  3.500 2.950 3.510 3.640 ;
        RECT  0.830 1.280 3.510 1.520 ;
        RECT  3.510 1.280 3.750 3.640 ;
        RECT  3.750 2.950 3.760 3.640 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.920 3.010 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 0.880 2.090 ;
        RECT  0.880 1.830 1.120 2.100 ;
        RECT  1.120 1.860 1.350 2.100 ;
        RECT  1.350 1.860 1.730 2.270 ;
        RECT  1.730 1.870 1.750 2.270 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.060 1.820 2.460 2.270 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.030 3.190 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.550 5.440 ;
        RECT  0.550 4.480 0.950 5.440 ;
        RECT  0.950 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.710 0.400 ;
        RECT  1.710 -0.400 2.110 0.560 ;
        RECT  2.110 -0.400 3.390 0.400 ;
        RECT  3.390 -0.400 3.790 0.560 ;
        RECT  3.790 -0.400 3.960 0.400 ;
        END
    END GND
END NOR4XL

MACRO NOR4X4
    CLASS CORE ;
    FOREIGN NOR4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR4XL ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.590 0.980 0.990 1.380 ;
        RECT  0.990 1.140 2.090 1.380 ;
        RECT  2.090 0.980 2.530 1.380 ;
        RECT  2.310 3.930 2.970 4.330 ;
        RECT  2.970 3.930 6.270 4.170 ;
        RECT  2.530 1.140 6.910 1.380 ;
        RECT  6.270 3.930 7.110 4.340 ;
        RECT  6.910 0.980 7.310 1.380 ;
        RECT  7.310 1.140 8.430 1.380 ;
        RECT  8.430 0.980 8.830 1.380 ;
        RECT  8.830 1.140 8.910 1.380 ;
        RECT  7.110 3.930 9.350 4.170 ;
        RECT  9.350 3.630 9.360 4.170 ;
        RECT  9.350 1.820 9.360 3.220 ;
        RECT  8.910 1.140 9.360 1.540 ;
        RECT  9.360 1.140 9.600 4.170 ;
        RECT  9.600 1.140 9.780 3.220 ;
        RECT  9.780 1.820 9.790 3.220 ;
        RECT  9.780 1.140 9.950 1.540 ;
        RECT  9.950 0.980 10.230 1.540 ;
        RECT  10.230 0.980 10.350 1.380 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.420 2.600 0.820 3.760 ;
        RECT  0.820 3.410 1.520 3.760 ;
        RECT  1.520 3.410 1.780 3.770 ;
        RECT  1.780 3.410 4.540 3.650 ;
        RECT  4.540 2.700 4.990 3.650 ;
        RECT  4.990 3.200 5.170 3.650 ;
        RECT  5.170 3.410 8.750 3.650 ;
        RECT  8.750 2.620 8.990 3.650 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 0.890 2.090 ;
        RECT  0.890 1.830 1.150 2.240 ;
        RECT  1.150 1.830 1.390 3.130 ;
        RECT  3.780 2.180 3.790 2.500 ;
        RECT  1.390 2.890 3.900 3.130 ;
        RECT  3.790 2.180 3.900 2.580 ;
        RECT  3.900 2.180 4.140 3.130 ;
        RECT  4.140 2.180 4.190 2.580 ;
        RECT  4.190 2.180 5.270 2.420 ;
        RECT  5.270 2.180 5.440 2.580 ;
        RECT  5.440 2.180 5.680 3.130 ;
        RECT  5.680 2.890 8.220 3.130 ;
        RECT  8.220 1.900 8.460 3.130 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.690 2.170 1.930 2.610 ;
        RECT  1.930 2.370 2.750 2.610 ;
        RECT  2.750 1.820 3.190 2.610 ;
        RECT  3.190 1.660 3.430 2.610 ;
        RECT  3.430 1.660 5.960 1.900 ;
        RECT  5.960 1.660 6.200 2.610 ;
        RECT  6.200 2.250 6.390 2.610 ;
        RECT  6.390 2.370 7.420 2.610 ;
        RECT  7.420 2.270 7.830 2.610 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.670 1.690 7.120 2.100 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.260 0.170 5.440 ;
        RECT  0.170 4.060 0.570 5.440 ;
        RECT  0.570 4.260 0.580 5.440 ;
        RECT  0.580 4.640 4.510 5.440 ;
        RECT  4.510 4.480 4.910 5.440 ;
        RECT  4.910 4.640 8.910 5.440 ;
        RECT  8.910 4.480 9.310 5.440 ;
        RECT  9.310 4.640 10.560 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.340 0.400 ;
        RECT  1.340 -0.400 1.350 0.740 ;
        RECT  1.350 -0.400 1.750 0.860 ;
        RECT  1.750 -0.400 1.760 0.740 ;
        RECT  1.760 -0.400 2.990 0.400 ;
        RECT  2.990 -0.400 3.000 0.740 ;
        RECT  3.000 -0.400 3.400 0.860 ;
        RECT  3.400 -0.400 3.410 0.740 ;
        RECT  3.410 -0.400 6.080 0.400 ;
        RECT  6.080 -0.400 6.090 0.740 ;
        RECT  6.090 -0.400 6.490 0.860 ;
        RECT  6.490 -0.400 6.500 0.740 ;
        RECT  6.500 -0.400 7.670 0.400 ;
        RECT  7.670 -0.400 8.070 0.850 ;
        RECT  8.070 -0.400 9.190 0.400 ;
        RECT  9.190 -0.400 9.590 0.850 ;
        RECT  9.590 -0.400 10.560 0.400 ;
        END
    END GND
END NOR4X4

MACRO NOR4X2
    CLASS CORE ;
    FOREIGN NOR4X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR4XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.950 4.130 4.410 4.370 ;
        RECT  4.410 4.080 4.510 4.370 ;
        RECT  4.510 4.060 4.670 4.370 ;
        RECT  1.170 0.860 4.820 1.100 ;
        RECT  4.670 3.940 4.910 4.370 ;
        RECT  4.820 0.710 5.080 1.100 ;
        RECT  5.080 0.860 5.390 1.100 ;
        RECT  4.910 3.940 5.550 4.180 ;
        RECT  5.390 0.860 5.550 1.280 ;
        RECT  5.550 0.860 5.790 4.180 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.780 2.400 0.860 2.800 ;
        RECT  0.860 2.390 1.120 2.800 ;
        RECT  1.120 2.400 1.180 2.800 ;
        RECT  1.180 2.560 2.090 2.800 ;
        RECT  2.090 2.560 2.350 2.960 ;
        RECT  2.350 2.560 2.590 3.750 ;
        RECT  2.590 3.500 2.750 3.750 ;
        RECT  2.750 3.510 4.120 3.750 ;
        RECT  4.120 3.420 4.360 3.750 ;
        RECT  4.360 3.420 4.730 3.660 ;
        RECT  4.730 3.200 5.020 3.660 ;
        RECT  5.020 2.410 5.260 3.660 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.500 1.860 1.520 2.260 ;
        RECT  1.520 1.830 1.660 2.260 ;
        RECT  1.660 1.380 1.900 2.260 ;
        RECT  1.900 1.380 4.620 1.620 ;
        RECT  4.620 1.380 4.860 2.050 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.230 1.970 4.050 2.210 ;
        RECT  4.050 1.970 4.290 2.650 ;
        RECT  4.290 2.390 4.420 2.650 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.990 2.500 3.320 2.740 ;
        RECT  3.320 2.500 3.500 3.200 ;
        RECT  3.500 2.500 3.560 3.210 ;
        RECT  3.560 2.950 3.760 3.210 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.750 5.440 ;
        RECT  0.750 3.130 1.150 5.440 ;
        RECT  1.150 4.640 5.300 5.440 ;
        RECT  5.300 4.480 5.700 5.440 ;
        RECT  5.700 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.350 0.400 ;
        RECT  0.350 -0.400 0.750 0.560 ;
        RECT  0.750 -0.400 1.990 0.400 ;
        RECT  1.990 -0.400 2.390 0.560 ;
        RECT  2.390 -0.400 3.700 0.400 ;
        RECT  3.700 -0.400 4.100 0.560 ;
        RECT  4.100 -0.400 5.940 0.400 ;
        END
    END GND
END NOR4X2

MACRO NOR4X1
    CLASS CORE ;
    FOREIGN NOR4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR4XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.930 1.150 1.330 1.550 ;
        RECT  1.330 1.260 1.530 1.550 ;
        RECT  1.530 1.310 2.430 1.550 ;
        RECT  2.430 1.260 2.570 1.550 ;
        RECT  2.570 1.150 2.970 1.550 ;
        RECT  2.750 3.360 3.060 3.760 ;
        RECT  3.060 3.360 3.410 3.770 ;
        RECT  3.410 3.220 3.510 3.770 ;
        RECT  2.970 1.310 3.510 1.550 ;
        RECT  3.510 1.310 3.750 3.770 ;
        RECT  3.750 3.510 3.760 3.770 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.610 3.000 ;
        RECT  0.610 2.420 1.000 3.000 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 0.880 2.090 ;
        RECT  0.880 1.830 0.980 2.100 ;
        RECT  0.980 1.830 1.120 2.180 ;
        RECT  1.120 1.860 1.350 2.180 ;
        RECT  1.350 1.860 1.750 2.260 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.050 1.820 2.450 2.270 ;
        RECT  2.450 1.820 2.520 2.100 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.760 2.390 3.140 2.970 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.540 5.440 ;
        RECT  0.540 4.480 0.940 5.440 ;
        RECT  0.940 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.750 0.400 ;
        RECT  1.750 -0.400 2.150 0.560 ;
        RECT  2.150 -0.400 3.390 0.400 ;
        RECT  3.390 -0.400 3.790 0.560 ;
        RECT  3.790 -0.400 3.960 0.400 ;
        END
    END GND
END NOR4X1

MACRO NOR3BXL
    CLASS CORE ;
    FOREIGN NOR3BXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.850 1.250 3.090 1.490 ;
        RECT  3.090 1.250 3.190 1.520 ;
        RECT  2.800 3.490 3.200 3.890 ;
        RECT  3.190 1.250 3.390 1.540 ;
        RECT  3.200 3.490 3.510 3.780 ;
        RECT  3.390 1.170 3.510 1.570 ;
        RECT  3.510 1.170 3.750 3.780 ;
        RECT  3.750 3.490 3.760 3.780 ;
        RECT  3.750 1.170 3.790 1.570 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.370 1.820 1.430 2.220 ;
        RECT  1.430 1.820 1.770 2.650 ;
        RECT  1.770 2.390 1.780 2.650 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.090 1.820 2.530 2.250 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.490 3.720 0.860 4.120 ;
        RECT  0.860 3.510 1.120 4.120 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.060 5.440 ;
        RECT  1.060 4.480 1.460 5.440 ;
        RECT  1.460 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.070 0.400 ;
        RECT  1.070 -0.400 1.470 0.560 ;
        RECT  1.470 -0.400 2.720 0.400 ;
        RECT  2.720 -0.400 3.120 0.560 ;
        RECT  3.120 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.790 2.530 2.950 2.930 ;
        RECT  2.550 2.530 2.790 3.180 ;
        RECT  0.490 2.940 2.550 3.180 ;
        RECT  0.490 1.310 0.580 1.710 ;
        RECT  0.250 1.310 0.490 3.450 ;
        RECT  0.180 1.310 0.250 1.710 ;
    END
END NOR3BXL

MACRO NOR3BX4
    CLASS CORE ;
    FOREIGN NOR3BX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR3BXL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.730 0.840 1.740 1.230 ;
        RECT  1.740 0.820 2.140 1.230 ;
        RECT  2.620 3.330 3.020 4.310 ;
        RECT  2.140 0.860 3.390 1.230 ;
        RECT  3.390 0.820 3.790 1.230 ;
        RECT  3.790 0.860 5.040 1.230 ;
        RECT  3.020 3.340 5.610 3.710 ;
        RECT  5.040 0.820 5.730 1.230 ;
        RECT  5.610 3.340 6.050 3.780 ;
        RECT  6.050 2.940 6.490 4.340 ;
        RECT  6.490 2.940 6.610 3.300 ;
        RECT  5.730 0.870 6.610 1.230 ;
        RECT  6.610 0.870 6.970 3.300 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.200 2.450 1.360 2.850 ;
        RECT  1.360 2.450 1.520 3.200 ;
        RECT  1.520 2.450 1.600 3.210 ;
        RECT  1.600 2.720 1.780 3.210 ;
        RECT  1.780 2.720 4.510 2.960 ;
        RECT  4.510 2.540 4.920 2.960 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.920 2.030 2.320 2.440 ;
        RECT  2.320 2.200 3.600 2.440 ;
        RECT  3.600 2.020 4.000 2.440 ;
        RECT  4.000 2.020 5.230 2.260 ;
        RECT  5.230 2.020 5.730 2.660 ;
        RECT  5.730 2.390 5.740 2.660 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 1.700 0.860 3.760 ;
        RECT  0.860 1.700 0.920 3.770 ;
        RECT  0.920 3.510 1.120 3.770 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.920 5.440 ;
        RECT  0.920 4.370 0.930 5.440 ;
        RECT  0.930 4.170 1.330 5.440 ;
        RECT  1.330 4.370 1.340 5.440 ;
        RECT  1.340 4.620 4.320 5.440 ;
        RECT  4.320 4.170 4.720 5.440 ;
        RECT  4.720 4.640 7.260 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.960 0.400 ;
        RECT  0.960 -0.400 0.970 0.700 ;
        RECT  0.970 -0.400 1.370 0.900 ;
        RECT  1.370 -0.400 1.380 0.700 ;
        RECT  1.380 -0.400 2.570 0.400 ;
        RECT  2.570 -0.400 2.970 0.560 ;
        RECT  2.970 -0.400 4.210 0.400 ;
        RECT  4.210 -0.400 4.610 0.560 ;
        RECT  4.610 -0.400 5.910 0.400 ;
        RECT  5.910 -0.400 6.310 0.560 ;
        RECT  6.310 -0.400 7.260 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.090 1.500 6.330 2.450 ;
        RECT  3.270 1.500 6.090 1.740 ;
        RECT  2.860 1.500 3.270 1.920 ;
        RECT  1.460 1.500 2.860 1.740 ;
        RECT  1.220 1.180 1.460 1.740 ;
        RECT  0.610 1.180 1.220 1.420 ;
        RECT  0.400 0.940 0.610 1.420 ;
        RECT  0.400 4.050 0.570 4.290 ;
        RECT  0.160 0.940 0.400 4.290 ;
    END
END NOR3BX4

MACRO NOR3BX2
    CLASS CORE ;
    FOREIGN NOR3BX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR3BXL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.870 0.800 1.930 1.200 ;
        RECT  1.930 0.800 2.270 1.210 ;
        RECT  2.620 3.460 3.020 3.860 ;
        RECT  2.270 0.860 3.530 1.210 ;
        RECT  3.530 0.800 4.170 1.210 ;
        RECT  3.020 3.500 4.650 3.780 ;
        RECT  4.170 0.930 4.650 1.210 ;
        RECT  4.650 0.930 4.930 3.780 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.160 2.420 1.520 2.660 ;
        RECT  1.520 2.390 1.540 2.660 ;
        RECT  1.540 1.480 1.780 2.660 ;
        RECT  1.780 1.480 1.870 1.820 ;
        RECT  1.870 1.480 4.130 1.720 ;
        RECT  4.130 1.480 4.370 2.640 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.140 2.010 2.380 2.620 ;
        RECT  2.380 2.010 2.430 2.400 ;
        RECT  2.430 2.010 2.530 2.380 ;
        RECT  2.530 2.010 3.410 2.250 ;
        RECT  3.410 2.010 3.730 2.650 ;
        RECT  3.730 2.390 3.760 2.650 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 1.620 0.770 2.020 ;
        RECT  0.770 1.270 1.120 2.020 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.920 5.440 ;
        RECT  0.920 3.920 0.930 5.440 ;
        RECT  0.930 3.720 1.330 5.440 ;
        RECT  1.330 3.920 1.340 5.440 ;
        RECT  1.340 4.640 4.390 5.440 ;
        RECT  4.390 4.480 4.790 5.440 ;
        RECT  4.790 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.040 0.400 ;
        RECT  1.040 -0.400 1.440 0.560 ;
        RECT  1.440 -0.400 2.700 0.400 ;
        RECT  2.700 -0.400 3.100 0.560 ;
        RECT  3.100 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.860 2.640 3.100 3.180 ;
        RECT  0.570 2.940 2.860 3.180 ;
        RECT  0.400 2.940 0.570 3.780 ;
        RECT  0.400 0.940 0.490 1.340 ;
        RECT  0.160 0.940 0.400 3.780 ;
    END
END NOR3BX2

MACRO NOR3BX1
    CLASS CORE ;
    FOREIGN NOR3BX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR3BXL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.720 0.970 3.410 1.210 ;
        RECT  2.880 3.610 3.510 4.010 ;
        RECT  3.500 1.830 3.510 2.090 ;
        RECT  3.410 0.970 3.510 1.500 ;
        RECT  3.510 0.970 3.750 4.010 ;
        RECT  3.750 1.830 3.760 2.090 ;
        RECT  3.750 0.970 3.780 1.500 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.470 2.240 1.830 2.810 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.980 1.550 2.180 1.950 ;
        RECT  2.180 1.550 2.430 2.090 ;
        RECT  2.430 1.830 2.440 2.090 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.740 1.780 1.140 2.270 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.120 5.440 ;
        RECT  1.120 4.480 1.520 5.440 ;
        RECT  1.520 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.890 0.400 ;
        RECT  0.890 -0.400 1.290 0.560 ;
        RECT  1.290 -0.400 2.560 0.400 ;
        RECT  2.560 -0.400 2.960 0.560 ;
        RECT  2.960 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.800 2.270 3.040 3.330 ;
        RECT  0.680 3.090 2.800 3.330 ;
        RECT  0.440 2.850 0.680 3.330 ;
        RECT  0.440 1.250 0.600 1.490 ;
        RECT  0.200 1.250 0.440 3.330 ;
    END
END NOR3BX1

MACRO NOR3XL
    CLASS CORE ;
    FOREIGN NOR3XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.180 1.160 0.580 1.560 ;
        RECT  0.580 1.260 0.770 1.560 ;
        RECT  0.770 1.280 0.870 1.560 ;
        RECT  0.870 1.320 1.770 1.560 ;
        RECT  1.770 1.280 1.870 1.560 ;
        RECT  1.870 1.160 2.270 1.560 ;
        RECT  1.920 3.180 2.320 3.580 ;
        RECT  2.320 3.180 2.850 3.420 ;
        RECT  2.270 1.270 2.850 1.560 ;
        RECT  2.850 1.270 3.090 3.420 ;
        RECT  3.090 1.270 3.100 1.560 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.190 2.390 0.890 2.980 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 1.120 2.090 ;
        RECT  1.120 1.840 1.620 2.080 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.390 1.670 2.650 ;
        RECT  1.670 2.390 2.070 2.880 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.180 5.440 ;
        RECT  0.180 4.480 0.580 5.440 ;
        RECT  0.580 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.060 0.400 ;
        RECT  1.060 -0.400 1.460 0.560 ;
        RECT  1.460 -0.400 2.740 0.400 ;
        RECT  2.740 -0.400 3.140 0.560 ;
        RECT  3.140 -0.400 3.300 0.400 ;
        END
    END GND
END NOR3XL

MACRO NOR3X4
    CLASS CORE ;
    FOREIGN NOR3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR3XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.920 0.800 0.930 1.210 ;
        RECT  0.930 0.780 1.330 1.210 ;
        RECT  2.050 3.660 2.540 4.080 ;
        RECT  1.330 0.850 2.570 1.210 ;
        RECT  2.570 0.780 2.970 1.210 ;
        RECT  2.970 0.850 4.210 1.210 ;
        RECT  4.210 0.780 4.610 1.210 ;
        RECT  2.540 3.660 4.820 3.900 ;
        RECT  4.820 3.470 5.390 3.900 ;
        RECT  5.390 2.380 5.650 3.900 ;
        RECT  5.650 2.380 5.890 4.060 ;
        RECT  4.610 0.850 5.890 1.210 ;
        RECT  5.890 0.850 6.050 4.060 ;
        RECT  6.050 0.850 6.250 3.220 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.410 1.690 0.860 3.210 ;
        RECT  0.860 2.950 1.120 3.210 ;
        RECT  1.120 2.960 3.620 3.200 ;
        RECT  3.620 2.940 3.960 3.200 ;
        RECT  3.960 2.600 4.360 3.200 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.260 1.650 1.500 2.610 ;
        RECT  1.500 2.370 2.840 2.610 ;
        RECT  2.840 2.370 3.030 2.650 ;
        RECT  3.030 2.080 3.100 2.650 ;
        RECT  3.100 2.080 3.430 2.610 ;
        RECT  3.430 2.080 4.770 2.320 ;
        RECT  4.770 2.080 5.010 2.890 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 1.830 2.260 2.090 ;
        RECT  2.260 1.480 2.670 2.090 ;
        RECT  2.670 1.480 5.380 1.720 ;
        RECT  5.380 1.480 5.620 1.880 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.230 5.440 ;
        RECT  0.230 4.070 0.240 5.440 ;
        RECT  0.240 3.580 0.640 5.440 ;
        RECT  0.640 4.070 0.650 5.440 ;
        RECT  0.650 4.610 3.720 5.440 ;
        RECT  3.720 4.360 3.730 5.440 ;
        RECT  3.730 4.240 4.130 5.440 ;
        RECT  4.130 4.360 4.140 5.440 ;
        RECT  4.140 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 0.930 ;
        RECT  0.170 -0.400 0.570 1.130 ;
        RECT  0.570 -0.400 0.580 0.930 ;
        RECT  0.580 -0.400 1.750 0.400 ;
        RECT  1.750 -0.400 2.150 0.560 ;
        RECT  2.150 -0.400 3.390 0.400 ;
        RECT  3.390 -0.400 3.790 0.560 ;
        RECT  3.790 -0.400 5.030 0.400 ;
        RECT  5.030 -0.400 5.430 0.560 ;
        RECT  5.430 -0.400 6.600 0.400 ;
        END
    END GND
END NOR3X4

MACRO NOR3X2
    CLASS CORE ;
    FOREIGN NOR3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR3XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.010 1.090 1.080 1.490 ;
        RECT  1.910 3.480 2.310 3.880 ;
        RECT  1.080 1.080 3.060 1.500 ;
        RECT  2.310 3.480 3.070 3.720 ;
        RECT  3.070 3.260 3.310 3.720 ;
        RECT  3.310 3.260 4.070 3.500 ;
        RECT  4.070 3.220 4.170 3.500 ;
        RECT  4.160 1.830 4.170 2.090 ;
        RECT  3.060 1.080 4.170 1.490 ;
        RECT  4.170 1.080 4.410 3.500 ;
        RECT  4.410 1.830 4.420 2.090 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.480 2.650 0.880 3.210 ;
        RECT  0.880 2.950 1.120 3.210 ;
        RECT  1.120 2.960 2.530 3.200 ;
        RECT  2.530 2.940 2.550 3.200 ;
        RECT  2.550 2.740 2.790 3.200 ;
        RECT  2.790 2.740 3.410 2.980 ;
        RECT  3.410 2.640 3.530 2.980 ;
        RECT  3.530 2.300 3.770 2.980 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.920 1.800 1.160 2.200 ;
        RECT  1.160 1.800 2.430 2.040 ;
        RECT  2.430 1.800 2.530 2.080 ;
        RECT  2.530 1.800 2.730 2.100 ;
        RECT  2.730 1.800 3.130 2.200 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.370 1.780 2.650 ;
        RECT  1.780 2.370 2.270 2.610 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.220 5.440 ;
        RECT  0.220 4.350 0.230 5.440 ;
        RECT  0.230 4.150 0.630 5.440 ;
        RECT  0.630 4.350 0.640 5.440 ;
        RECT  0.640 4.640 3.580 5.440 ;
        RECT  3.580 4.000 3.590 5.440 ;
        RECT  3.590 3.800 3.990 5.440 ;
        RECT  3.990 4.000 4.000 5.440 ;
        RECT  4.000 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.760 0.400 ;
        RECT  1.760 -0.400 1.770 0.690 ;
        RECT  1.770 -0.400 2.170 0.810 ;
        RECT  2.170 -0.400 2.180 0.690 ;
        RECT  2.180 -0.400 3.740 0.400 ;
        RECT  3.740 -0.400 3.750 0.680 ;
        RECT  3.750 -0.400 4.150 0.800 ;
        RECT  4.150 -0.400 4.160 0.680 ;
        RECT  4.160 -0.400 4.620 0.400 ;
        END
    END GND
END NOR3X2

MACRO NOR3X1
    CLASS CORE ;
    FOREIGN NOR3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR3XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.990 1.150 1.390 1.550 ;
        RECT  1.390 1.260 1.530 1.550 ;
        RECT  1.920 3.510 2.320 3.910 ;
        RECT  1.530 1.310 2.430 1.550 ;
        RECT  2.320 3.510 2.530 3.780 ;
        RECT  2.430 1.260 2.630 1.550 ;
        RECT  2.530 3.500 2.750 3.780 ;
        RECT  2.630 1.220 2.750 1.620 ;
        RECT  2.750 1.220 2.990 3.780 ;
        RECT  2.990 1.220 3.030 1.840 ;
        RECT  2.990 3.510 3.100 3.780 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.460 3.030 ;
        RECT  0.460 2.630 0.880 3.030 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 1.120 2.180 ;
        RECT  1.120 1.940 1.590 2.180 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.950 1.670 3.210 ;
        RECT  1.670 2.640 2.070 3.210 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.220 0.400 ;
        RECT  0.220 -0.400 0.640 1.560 ;
        RECT  0.640 -0.400 1.810 0.400 ;
        RECT  1.810 -0.400 2.210 0.560 ;
        RECT  2.210 -0.400 3.300 0.400 ;
        END
    END GND
END NOR3X1

MACRO NOR2BXL
    CLASS CORE ;
    FOREIGN NOR2BXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.450 1.280 2.850 1.680 ;
        RECT  2.790 3.510 2.890 4.100 ;
        RECT  2.850 1.440 2.890 1.840 ;
        RECT  2.890 1.440 3.130 4.100 ;
        RECT  3.130 3.510 3.140 4.100 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.490 2.650 1.880 3.220 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.850 1.820 1.220 2.420 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.440 5.440 ;
        RECT  1.440 4.480 1.840 5.440 ;
        RECT  1.840 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.270 0.400 ;
        RECT  1.270 -0.400 1.670 0.560 ;
        RECT  1.670 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.470 2.250 2.610 2.650 ;
        RECT  2.230 1.970 2.470 3.720 ;
        RECT  2.180 1.970 2.230 2.210 ;
        RECT  0.930 3.480 2.230 3.720 ;
        RECT  1.940 1.300 2.180 2.210 ;
        RECT  0.390 1.300 1.940 1.540 ;
        RECT  0.530 3.480 0.930 3.880 ;
    END
END NOR2BXL

MACRO NOR2BX4
    CLASS CORE ;
    FOREIGN NOR2BX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR2BXL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.690 0.930 2.090 1.440 ;
        RECT  2.090 1.080 3.210 1.440 ;
        RECT  3.210 0.930 3.610 1.440 ;
        RECT  2.260 2.910 4.070 3.330 ;
        RECT  4.070 2.910 4.510 4.340 ;
        RECT  4.510 2.910 4.670 3.260 ;
        RECT  4.670 2.850 4.730 3.260 ;
        RECT  4.730 2.520 4.760 3.260 ;
        RECT  3.610 1.080 4.760 1.440 ;
        RECT  4.760 1.080 5.120 3.260 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.450 1.770 1.850 2.120 ;
        RECT  1.850 1.770 3.440 2.010 ;
        RECT  3.440 1.770 3.840 2.120 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.130 1.830 0.500 2.420 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.880 5.440 ;
        RECT  0.880 4.160 0.890 5.440 ;
        RECT  0.890 4.040 1.290 5.440 ;
        RECT  1.290 4.160 1.300 5.440 ;
        RECT  1.300 4.640 3.400 5.440 ;
        RECT  3.400 3.850 3.800 5.440 ;
        RECT  3.800 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.920 0.400 ;
        RECT  0.920 -0.400 0.930 0.710 ;
        RECT  0.930 -0.400 1.330 0.910 ;
        RECT  1.330 -0.400 1.340 0.710 ;
        RECT  1.340 -0.400 2.440 0.400 ;
        RECT  2.440 -0.400 2.450 0.690 ;
        RECT  2.450 -0.400 2.850 0.810 ;
        RECT  2.850 -0.400 2.860 0.690 ;
        RECT  2.860 -0.400 4.010 0.400 ;
        RECT  4.010 -0.400 4.410 0.560 ;
        RECT  4.410 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.240 1.800 4.480 2.640 ;
        RECT  2.620 2.400 4.240 2.640 ;
        RECT  2.220 2.320 2.620 2.640 ;
        RECT  1.050 2.400 2.220 2.640 ;
        RECT  0.810 1.230 1.050 3.740 ;
        RECT  0.570 1.230 0.810 1.550 ;
        RECT  0.170 3.500 0.810 3.740 ;
        RECT  0.170 1.150 0.570 1.550 ;
    END
END NOR2BX4

MACRO NOR2BX2
    CLASS CORE ;
    FOREIGN NOR2BX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR2BXL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.670 0.820 2.070 1.220 ;
        RECT  2.280 3.660 2.840 3.900 ;
        RECT  2.840 3.510 3.100 3.900 ;
        RECT  2.070 0.980 3.410 1.220 ;
        RECT  3.100 3.660 3.480 3.900 ;
        RECT  3.410 0.980 3.480 1.260 ;
        RECT  3.480 0.980 3.720 3.900 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.300 2.550 1.520 2.790 ;
        RECT  1.520 1.790 1.780 2.790 ;
        RECT  1.780 1.790 2.960 2.070 ;
        RECT  2.960 1.790 2.970 2.200 ;
        RECT  2.970 1.800 3.200 2.200 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 1.750 0.770 2.170 ;
        RECT  0.770 1.270 1.110 2.170 ;
        RECT  1.110 1.270 1.120 1.530 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.970 5.440 ;
        RECT  0.970 3.710 0.980 5.440 ;
        RECT  0.980 3.590 1.380 5.440 ;
        RECT  1.380 3.710 1.390 5.440 ;
        RECT  1.390 4.640 3.400 5.440 ;
        RECT  3.400 4.480 3.800 5.440 ;
        RECT  3.800 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.860 0.400 ;
        RECT  0.860 -0.400 1.260 0.560 ;
        RECT  1.260 -0.400 2.480 0.400 ;
        RECT  2.480 -0.400 2.880 0.560 ;
        RECT  2.880 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.400 2.350 2.570 2.590 ;
        RECT  2.160 2.350 2.400 3.310 ;
        RECT  0.570 3.070 2.160 3.310 ;
        RECT  0.400 3.070 0.570 3.510 ;
        RECT  0.400 1.060 0.490 1.460 ;
        RECT  0.160 1.060 0.400 3.510 ;
    END
END NOR2BX2

MACRO NOR2BX1
    CLASS CORE ;
    FOREIGN NOR2BX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR2BXL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.720 0.950 2.120 1.350 ;
        RECT  2.420 3.060 2.760 4.040 ;
        RECT  2.120 1.110 2.760 1.350 ;
        RECT  2.760 1.110 2.820 4.040 ;
        RECT  2.820 1.110 3.000 3.310 ;
        RECT  3.000 1.830 3.100 2.090 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 1.700 2.000 2.100 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.720 2.340 1.210 2.740 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.120 5.440 ;
        RECT  1.120 4.480 1.520 5.440 ;
        RECT  1.520 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.890 0.400 ;
        RECT  0.890 -0.400 1.290 0.560 ;
        RECT  1.290 -0.400 2.580 0.400 ;
        RECT  2.580 -0.400 2.980 0.560 ;
        RECT  2.980 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.140 2.390 2.480 2.790 ;
        RECT  1.900 2.390 2.140 3.450 ;
        RECT  0.600 3.210 1.900 3.450 ;
        RECT  0.440 1.170 0.600 1.570 ;
        RECT  0.440 3.020 0.600 3.450 ;
        RECT  0.200 1.170 0.440 3.450 ;
    END
END NOR2BX1

MACRO NOR2XL
    CLASS CORE ;
    FOREIGN NOR2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 3.510 1.530 3.770 ;
        RECT  1.530 2.940 1.780 3.770 ;
        RECT  1.010 1.280 1.870 1.520 ;
        RECT  1.780 2.940 1.980 3.680 ;
        RECT  1.870 1.280 1.980 1.540 ;
        RECT  1.980 1.280 2.020 3.680 ;
        RECT  2.020 1.280 2.220 3.180 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.190 2.390 0.950 2.980 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 1.120 2.090 ;
        RECT  1.120 1.840 1.460 2.080 ;
        RECT  1.460 1.840 1.700 2.360 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.360 5.440 ;
        RECT  0.360 4.480 0.760 5.440 ;
        RECT  0.760 4.640 2.640 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.190 0.400 ;
        RECT  0.190 -0.400 0.590 0.560 ;
        RECT  0.590 -0.400 1.890 0.400 ;
        RECT  1.890 -0.400 2.290 0.560 ;
        RECT  2.290 -0.400 2.640 0.400 ;
        END
    END GND
END NOR2XL

MACRO NOR2X4
    CLASS CORE ;
    FOREIGN NOR2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR2XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.890 1.030 1.290 1.430 ;
        RECT  1.290 1.190 2.330 1.430 ;
        RECT  2.330 1.030 2.350 1.430 ;
        RECT  2.350 1.030 2.730 1.440 ;
        RECT  1.530 2.920 4.070 3.320 ;
        RECT  4.070 2.380 4.140 3.780 ;
        RECT  2.730 1.080 4.140 1.440 ;
        RECT  4.140 1.080 4.500 3.780 ;
        RECT  4.500 2.380 4.760 3.780 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.460 2.250 0.860 2.650 ;
        RECT  0.860 2.390 1.120 2.650 ;
        RECT  1.120 2.400 2.430 2.640 ;
        RECT  2.430 2.330 3.140 2.640 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.530 2.090 ;
        RECT  1.530 1.760 1.690 2.090 ;
        RECT  1.690 1.760 2.190 2.120 ;
        RECT  2.190 1.760 3.490 2.000 ;
        RECT  3.490 1.760 3.890 2.110 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 3.060 5.440 ;
        RECT  3.060 3.850 3.460 5.440 ;
        RECT  3.460 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 0.710 ;
        RECT  0.170 -0.400 0.570 0.910 ;
        RECT  0.570 -0.400 0.580 0.710 ;
        RECT  0.580 -0.400 1.600 0.400 ;
        RECT  1.600 -0.400 2.020 0.920 ;
        RECT  2.020 -0.400 3.130 0.400 ;
        RECT  3.130 -0.400 3.530 0.560 ;
        RECT  3.530 -0.400 5.280 0.400 ;
        END
    END GND
END NOR2X4

MACRO NOR2X2
    CLASS CORE ;
    FOREIGN NOR2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR2XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.130 1.090 1.330 1.490 ;
        RECT  1.430 3.030 1.830 3.430 ;
        RECT  1.830 3.030 2.850 3.270 ;
        RECT  2.840 2.390 2.850 2.650 ;
        RECT  1.330 1.080 2.850 1.500 ;
        RECT  2.850 1.080 2.930 3.270 ;
        RECT  2.930 1.090 3.090 3.270 ;
        RECT  3.090 2.390 3.100 2.650 ;
        RECT  3.090 1.090 3.130 1.490 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.490 1.800 0.890 2.630 ;
        RECT  0.890 1.800 1.120 2.090 ;
        RECT  1.120 1.800 2.240 2.040 ;
        RECT  2.240 1.800 2.480 2.200 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.300 2.360 1.870 2.740 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 2.690 5.440 ;
        RECT  2.690 4.480 3.090 5.440 ;
        RECT  3.090 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.930 0.400 ;
        RECT  1.930 -0.400 2.330 0.560 ;
        RECT  2.330 -0.400 3.300 0.400 ;
        END
    END GND
END NOR2X2

MACRO NOR2X1
    CLASS CORE ;
    FOREIGN NOR2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NOR2XL ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.750 1.150 1.150 1.550 ;
        RECT  1.410 3.230 1.430 3.640 ;
        RECT  1.430 3.220 1.490 3.640 ;
        RECT  1.490 2.920 1.580 3.640 ;
        RECT  1.150 1.310 1.580 1.550 ;
        RECT  1.580 1.310 1.820 3.640 ;
        RECT  1.820 3.050 1.830 3.640 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.150 2.260 0.500 2.980 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 1.300 2.260 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.980 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.400 0.400 ;
        RECT  1.400 -0.400 1.800 0.560 ;
        RECT  1.800 -0.400 1.980 0.400 ;
        END
    END GND
END NOR2X1

MACRO NAND4BBXL
    CLASS CORE ;
    FOREIGN NAND4BBXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.730 3.520 2.130 3.920 ;
        RECT  2.130 3.520 3.190 3.760 ;
        RECT  3.190 3.520 3.230 3.780 ;
        RECT  3.230 3.520 3.500 3.920 ;
        RECT  3.500 3.510 3.630 3.920 ;
        RECT  3.630 3.510 3.760 3.770 ;
        RECT  3.520 1.320 3.760 2.610 ;
        RECT  3.760 3.520 4.200 3.760 ;
        RECT  3.760 2.370 4.200 2.610 ;
        RECT  4.200 2.370 4.440 3.760 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.360 2.040 1.370 2.580 ;
        RECT  1.370 1.840 1.520 2.580 ;
        RECT  1.520 1.830 1.620 2.580 ;
        RECT  1.620 1.830 1.780 2.090 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.000 2.380 2.530 2.720 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.030 1.680 4.510 2.100 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.020 0.580 3.020 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.040 5.440 ;
        RECT  1.040 4.480 1.440 5.440 ;
        RECT  1.440 4.640 2.420 5.440 ;
        RECT  2.420 4.480 2.820 5.440 ;
        RECT  2.820 4.640 3.940 5.440 ;
        RECT  3.940 4.480 4.340 5.440 ;
        RECT  4.340 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.240 0.400 ;
        RECT  1.240 -0.400 1.640 0.560 ;
        RECT  1.640 -0.400 4.630 0.400 ;
        RECT  4.630 -0.400 5.030 0.560 ;
        RECT  5.030 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.790 1.170 5.030 3.750 ;
        RECT  4.280 1.170 4.790 1.410 ;
        RECT  4.040 0.750 4.280 1.410 ;
        RECT  3.240 0.750 4.040 0.990 ;
        RECT  3.520 2.890 3.920 3.230 ;
        RECT  1.090 2.990 3.520 3.230 ;
        RECT  3.000 0.750 3.240 2.640 ;
        RECT  2.800 2.400 3.000 2.640 ;
        RECT  0.850 1.310 1.090 3.730 ;
        RECT  0.760 1.310 0.850 1.550 ;
        RECT  0.570 3.490 0.850 3.730 ;
        RECT  0.360 1.150 0.760 1.550 ;
        RECT  0.170 3.490 0.570 3.890 ;
    END
END NAND4BBXL

MACRO NAND4BBX4
    CLASS CORE ;
    FOREIGN NAND4BBX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND4BBXL ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 3.660 2.580 4.060 ;
        RECT  2.580 3.660 3.820 3.900 ;
        RECT  3.820 3.660 4.220 4.060 ;
        RECT  3.850 0.670 5.530 0.910 ;
        RECT  5.530 0.670 5.770 1.100 ;
        RECT  4.220 3.660 8.490 3.900 ;
        RECT  8.490 3.660 8.890 4.060 ;
        RECT  8.890 3.660 9.570 3.900 ;
        RECT  9.570 3.500 10.010 3.900 ;
        RECT  10.010 2.940 10.450 4.340 ;
        RECT  10.450 3.500 10.530 4.060 ;
        RECT  10.530 3.500 10.890 3.900 ;
        RECT  5.770 0.860 12.650 1.100 ;
        RECT  10.890 3.660 12.700 3.900 ;
        RECT  12.650 0.860 12.700 1.400 ;
        RECT  12.700 0.860 12.940 3.900 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.390 1.190 1.630 2.240 ;
        RECT  1.630 1.190 4.820 1.430 ;
        RECT  4.820 1.190 5.080 1.620 ;
        RECT  5.080 1.380 6.050 1.620 ;
        RECT  6.050 1.380 6.490 1.940 ;
        RECT  6.490 1.380 10.880 1.620 ;
        RECT  10.880 1.380 11.120 2.150 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.430 2.300 2.590 2.540 ;
        RECT  2.590 2.300 2.880 3.320 ;
        RECT  2.880 3.080 5.630 3.320 ;
        RECT  5.630 2.980 6.030 3.380 ;
        RECT  6.030 2.980 6.810 3.220 ;
        RECT  6.810 2.980 7.210 3.380 ;
        RECT  7.210 2.980 8.120 3.220 ;
        RECT  8.120 2.950 8.380 3.220 ;
        RECT  8.380 2.960 9.500 3.220 ;
        RECT  9.500 2.420 9.740 3.220 ;
        RECT  9.740 2.420 10.070 2.660 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  11.920 2.080 12.340 2.650 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.020 0.590 2.650 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.260 5.440 ;
        RECT  1.260 4.480 1.660 5.440 ;
        RECT  1.660 4.640 3.000 5.440 ;
        RECT  3.000 4.480 3.400 5.440 ;
        RECT  3.400 4.640 4.570 5.440 ;
        RECT  4.570 4.300 4.580 5.440 ;
        RECT  4.580 4.180 4.980 5.440 ;
        RECT  4.980 4.300 4.990 5.440 ;
        RECT  4.990 4.640 7.720 5.440 ;
        RECT  7.720 4.300 7.730 5.440 ;
        RECT  7.730 4.180 8.130 5.440 ;
        RECT  8.130 4.300 8.140 5.440 ;
        RECT  8.140 4.640 9.310 5.440 ;
        RECT  9.310 4.480 9.710 5.440 ;
        RECT  9.710 4.640 10.950 5.440 ;
        RECT  10.950 4.480 11.350 5.440 ;
        RECT  11.350 4.640 13.200 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.120 0.400 ;
        RECT  1.120 -0.400 2.100 0.910 ;
        RECT  2.100 -0.400 6.050 0.400 ;
        RECT  6.050 -0.400 6.450 0.560 ;
        RECT  6.450 -0.400 10.470 0.400 ;
        RECT  10.470 -0.400 11.450 0.560 ;
        RECT  11.450 -0.400 13.200 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  11.640 1.380 12.390 1.620 ;
        RECT  11.640 2.930 12.170 3.330 ;
        RECT  11.400 1.380 11.640 3.330 ;
        RECT  10.590 2.430 11.400 2.670 ;
        RECT  10.350 1.900 10.590 2.670 ;
        RECT  9.010 1.900 10.350 2.140 ;
        RECT  8.770 1.900 9.010 2.660 ;
        RECT  7.930 2.420 8.770 2.660 ;
        RECT  7.530 2.130 7.930 2.660 ;
        RECT  5.310 2.420 7.530 2.660 ;
        RECT  4.910 2.420 5.310 2.800 ;
        RECT  3.710 2.420 4.910 2.660 ;
        RECT  2.150 1.740 4.470 1.980 ;
        RECT  3.290 2.280 3.710 2.660 ;
        RECT  1.910 1.740 2.150 2.760 ;
        RECT  1.110 2.520 1.910 2.760 ;
        RECT  0.870 1.310 1.110 3.730 ;
        RECT  0.740 1.310 0.870 1.550 ;
        RECT  0.750 3.490 0.870 3.730 ;
        RECT  0.350 3.490 0.750 4.370 ;
        RECT  0.340 0.670 0.740 1.550 ;
    END
END NAND4BBX4

MACRO NAND4BBX2
    CLASS CORE ;
    FOREIGN NAND4BBX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND4BBXL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.750 0.860 4.820 1.100 ;
        RECT  4.820 0.710 5.080 1.100 ;
        RECT  1.860 3.870 7.370 4.110 ;
        RECT  7.370 3.780 7.460 4.110 ;
        RECT  5.080 0.860 7.460 1.100 ;
        RECT  7.460 0.860 7.700 4.110 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.390 1.580 2.650 ;
        RECT  1.580 2.240 1.820 3.510 ;
        RECT  1.820 3.220 1.870 3.510 ;
        RECT  1.870 3.270 5.450 3.510 ;
        RECT  5.450 3.270 5.850 3.580 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 1.830 2.380 2.090 ;
        RECT  2.380 1.830 2.440 2.990 ;
        RECT  2.440 1.840 2.620 2.990 ;
        RECT  2.620 2.750 5.190 2.990 ;
        RECT  5.190 2.610 5.590 2.990 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.720 2.060 6.800 2.460 ;
        RECT  6.800 2.060 7.050 2.650 ;
        RECT  7.050 2.390 7.060 2.650 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.770 1.820 1.170 2.270 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.040 5.440 ;
        RECT  1.040 4.480 1.440 5.440 ;
        RECT  1.440 4.640 2.410 5.440 ;
        RECT  2.410 4.450 2.880 5.440 ;
        RECT  2.880 4.480 3.080 5.440 ;
        RECT  3.080 4.640 4.330 5.440 ;
        RECT  4.330 4.480 4.730 5.440 ;
        RECT  4.730 4.640 6.960 5.440 ;
        RECT  6.960 4.480 7.360 5.440 ;
        RECT  7.360 4.640 7.920 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.550 0.400 ;
        RECT  1.550 -0.400 1.950 0.560 ;
        RECT  1.950 -0.400 5.980 0.400 ;
        RECT  5.980 -0.400 6.380 0.560 ;
        RECT  6.380 -0.400 7.920 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.940 1.380 7.180 1.780 ;
        RECT  6.440 1.540 6.940 1.780 ;
        RECT  6.440 3.120 6.610 3.520 ;
        RECT  6.200 1.540 6.440 3.520 ;
        RECT  4.870 2.090 6.200 2.330 ;
        RECT  4.470 2.050 4.870 2.460 ;
        RECT  3.430 2.220 4.470 2.460 ;
        RECT  3.750 1.630 4.150 1.940 ;
        RECT  3.470 1.630 3.750 1.870 ;
        RECT  3.230 1.310 3.470 1.870 ;
        RECT  3.030 2.150 3.430 2.460 ;
        RECT  1.130 1.310 3.230 1.550 ;
        RECT  0.730 1.060 1.130 1.550 ;
        RECT  0.490 1.310 0.730 1.550 ;
        RECT  0.490 2.800 0.570 3.200 ;
        RECT  0.250 1.310 0.490 3.200 ;
        RECT  0.170 2.800 0.250 3.200 ;
    END
END NAND4BBX2

MACRO NAND4BBX1
    CLASS CORE ;
    FOREIGN NAND4BBX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND4BBXL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.730 3.520 2.130 3.920 ;
        RECT  2.130 3.520 3.190 3.760 ;
        RECT  3.190 3.520 3.230 3.780 ;
        RECT  3.230 3.520 3.500 3.920 ;
        RECT  3.500 3.510 3.630 3.920 ;
        RECT  3.630 3.510 3.760 3.770 ;
        RECT  3.520 1.320 3.760 2.610 ;
        RECT  3.760 3.510 4.200 3.760 ;
        RECT  3.760 2.370 4.200 2.610 ;
        RECT  4.200 2.370 4.440 3.760 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.360 1.830 1.620 2.700 ;
        RECT  1.620 1.830 1.780 2.090 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.000 2.380 2.530 2.720 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.030 1.680 4.510 2.100 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.820 0.580 2.650 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.040 5.440 ;
        RECT  1.040 4.480 1.440 5.440 ;
        RECT  1.440 4.640 2.420 5.440 ;
        RECT  2.420 4.480 2.820 5.440 ;
        RECT  2.820 4.640 4.040 5.440 ;
        RECT  4.040 4.480 4.440 5.440 ;
        RECT  4.440 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.240 0.400 ;
        RECT  1.240 -0.400 1.640 0.560 ;
        RECT  1.640 -0.400 4.710 0.400 ;
        RECT  4.710 -0.400 5.110 0.560 ;
        RECT  5.110 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.780 1.170 5.020 3.770 ;
        RECT  4.280 1.170 4.780 1.410 ;
        RECT  4.040 0.800 4.280 1.410 ;
        RECT  3.240 0.800 4.040 1.040 ;
        RECT  3.520 2.890 3.920 3.230 ;
        RECT  1.090 2.990 3.520 3.230 ;
        RECT  3.000 0.800 3.240 2.710 ;
        RECT  2.800 2.470 3.000 2.710 ;
        RECT  0.850 1.310 1.090 3.720 ;
        RECT  0.760 1.310 0.850 1.550 ;
        RECT  0.570 3.480 0.850 3.720 ;
        RECT  0.360 1.150 0.760 1.550 ;
        RECT  0.170 3.480 0.570 3.880 ;
    END
END NAND4BBX1

MACRO NAND4BXL
    CLASS CORE ;
    FOREIGN NAND4BXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.730 3.000 2.130 3.400 ;
        RECT  2.130 3.000 3.230 3.240 ;
        RECT  3.230 3.000 3.630 3.400 ;
        RECT  3.440 0.920 3.650 1.320 ;
        RECT  3.650 0.910 4.160 1.320 ;
        RECT  3.630 3.000 4.170 3.240 ;
        RECT  4.160 0.910 4.170 1.530 ;
        RECT  4.170 0.910 4.410 3.240 ;
        RECT  4.410 0.910 4.420 1.530 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 1.600 1.880 2.100 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.940 2.380 2.530 2.680 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.800 2.320 3.200 2.720 ;
        RECT  3.200 2.380 3.770 2.660 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.740 1.800 0.770 2.200 ;
        RECT  0.770 1.800 0.820 2.620 ;
        RECT  0.820 1.800 1.140 2.660 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.040 5.440 ;
        RECT  1.040 4.480 1.440 5.440 ;
        RECT  1.440 4.640 2.420 5.440 ;
        RECT  2.420 4.480 2.820 5.440 ;
        RECT  2.820 4.640 3.940 5.440 ;
        RECT  3.940 4.480 4.340 5.440 ;
        RECT  4.340 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.240 0.400 ;
        RECT  1.240 -0.400 1.640 0.560 ;
        RECT  1.640 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.200 1.600 3.600 2.000 ;
        RECT  3.160 1.600 3.200 1.840 ;
        RECT  2.920 1.080 3.160 1.840 ;
        RECT  0.760 1.080 2.920 1.320 ;
        RECT  0.480 1.080 0.760 1.550 ;
        RECT  0.480 2.900 0.570 3.300 ;
        RECT  0.240 1.080 0.480 3.300 ;
        RECT  0.170 2.900 0.240 3.300 ;
    END
END NAND4BXL

MACRO NAND4BX4
    CLASS CORE ;
    FOREIGN NAND4BX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND4BXL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 3.660 2.580 4.060 ;
        RECT  2.580 3.660 3.820 3.900 ;
        RECT  3.820 3.660 4.220 4.060 ;
        RECT  3.850 0.670 5.530 0.910 ;
        RECT  5.530 0.670 5.770 1.100 ;
        RECT  4.220 3.660 8.490 3.900 ;
        RECT  8.490 3.660 8.890 4.060 ;
        RECT  8.890 3.660 9.560 3.900 ;
        RECT  9.560 3.500 10.010 3.900 ;
        RECT  10.010 2.940 10.450 4.340 ;
        RECT  10.450 3.660 10.530 4.060 ;
        RECT  10.450 2.940 11.140 3.220 ;
        RECT  5.770 0.860 11.140 1.100 ;
        RECT  11.140 0.860 11.380 3.220 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.470 1.190 1.710 2.240 ;
        RECT  1.710 1.190 4.820 1.430 ;
        RECT  4.820 1.190 4.830 1.530 ;
        RECT  4.830 1.190 5.070 1.620 ;
        RECT  5.070 1.270 5.080 1.620 ;
        RECT  5.080 1.380 6.050 1.620 ;
        RECT  6.050 1.380 6.490 1.940 ;
        RECT  6.490 1.380 10.540 1.620 ;
        RECT  10.540 1.380 10.780 2.130 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.510 2.280 2.910 3.320 ;
        RECT  2.910 3.080 5.630 3.320 ;
        RECT  5.630 2.950 6.030 3.380 ;
        RECT  6.030 2.950 6.820 3.220 ;
        RECT  6.820 2.950 7.590 3.380 ;
        RECT  7.590 2.950 8.380 3.210 ;
        RECT  8.380 2.950 9.500 3.200 ;
        RECT  9.500 2.360 9.740 3.200 ;
        RECT  9.740 2.360 10.140 2.600 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.220 2.260 3.460 2.660 ;
        RECT  3.460 2.390 3.760 2.660 ;
        RECT  3.760 2.420 4.910 2.660 ;
        RECT  4.910 2.420 5.310 2.800 ;
        RECT  5.310 2.420 7.530 2.660 ;
        RECT  7.530 2.130 7.950 2.660 ;
        RECT  7.950 2.380 8.250 2.660 ;
        RECT  8.250 2.420 8.820 2.660 ;
        RECT  8.820 2.260 9.220 2.660 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.020 0.670 2.650 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.310 5.440 ;
        RECT  1.310 4.480 1.710 5.440 ;
        RECT  1.710 4.640 3.000 5.440 ;
        RECT  3.000 4.480 3.400 5.440 ;
        RECT  3.400 4.640 4.570 5.440 ;
        RECT  4.570 4.300 4.580 5.440 ;
        RECT  4.580 4.180 4.980 5.440 ;
        RECT  4.980 4.300 4.990 5.440 ;
        RECT  4.990 4.640 7.720 5.440 ;
        RECT  7.720 4.300 7.730 5.440 ;
        RECT  7.730 4.180 8.130 5.440 ;
        RECT  8.130 4.300 8.140 5.440 ;
        RECT  8.140 4.640 9.310 5.440 ;
        RECT  9.310 4.480 9.710 5.440 ;
        RECT  9.710 4.640 10.950 5.440 ;
        RECT  10.950 3.820 11.350 5.440 ;
        RECT  11.350 4.640 11.880 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.140 0.400 ;
        RECT  1.140 -0.400 2.120 0.910 ;
        RECT  2.120 -0.400 6.050 0.400 ;
        RECT  6.050 -0.400 6.450 0.560 ;
        RECT  6.450 -0.400 10.410 0.400 ;
        RECT  10.410 -0.400 10.810 0.560 ;
        RECT  10.810 -0.400 11.880 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.230 1.740 4.400 1.980 ;
        RECT  1.990 1.740 2.230 2.760 ;
        RECT  1.190 2.520 1.990 2.760 ;
        RECT  0.950 1.310 1.190 3.730 ;
        RECT  0.790 1.310 0.950 1.550 ;
        RECT  0.830 3.490 0.950 3.730 ;
        RECT  0.430 3.490 0.830 4.370 ;
        RECT  0.780 0.790 0.790 1.550 ;
        RECT  0.380 0.670 0.780 1.550 ;
        RECT  0.370 0.790 0.380 1.350 ;
    END
END NAND4BX4

MACRO NAND4BX2
    CLASS CORE ;
    FOREIGN NAND4BX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND4BXL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.750 0.790 5.390 1.030 ;
        RECT  5.390 0.790 5.630 1.530 ;
        RECT  1.860 3.870 6.130 4.110 ;
        RECT  5.630 1.260 6.130 1.530 ;
        RECT  6.130 1.260 6.370 4.110 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.390 1.580 2.650 ;
        RECT  1.580 2.240 1.820 3.510 ;
        RECT  1.820 3.220 1.870 3.510 ;
        RECT  1.870 3.270 5.450 3.510 ;
        RECT  5.450 3.270 5.850 3.580 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 1.830 2.380 2.090 ;
        RECT  2.380 1.830 2.440 2.990 ;
        RECT  2.440 1.840 2.620 2.990 ;
        RECT  2.620 2.750 5.180 2.990 ;
        RECT  5.180 2.530 5.580 2.990 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.030 2.070 3.430 2.470 ;
        RECT  3.430 2.220 4.470 2.460 ;
        RECT  4.470 2.050 4.630 2.460 ;
        RECT  4.630 1.840 4.820 2.460 ;
        RECT  4.820 1.830 4.870 2.460 ;
        RECT  4.870 1.830 5.080 2.090 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.770 1.820 1.170 2.270 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.040 5.440 ;
        RECT  1.040 4.480 1.440 5.440 ;
        RECT  1.440 4.640 2.680 5.440 ;
        RECT  2.680 4.480 3.080 5.440 ;
        RECT  3.080 4.640 4.330 5.440 ;
        RECT  4.330 4.480 4.730 5.440 ;
        RECT  4.730 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.550 0.400 ;
        RECT  1.550 -0.400 1.950 0.560 ;
        RECT  1.950 -0.400 5.980 0.400 ;
        RECT  5.980 -0.400 6.380 0.560 ;
        RECT  6.380 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.990 1.700 4.150 1.940 ;
        RECT  3.750 1.310 3.990 1.940 ;
        RECT  1.130 1.310 3.750 1.550 ;
        RECT  0.730 1.060 1.130 1.550 ;
        RECT  0.490 1.310 0.730 1.550 ;
        RECT  0.490 2.800 0.570 3.200 ;
        RECT  0.250 1.310 0.490 3.200 ;
        RECT  0.170 2.800 0.250 3.200 ;
    END
END NAND4BX2

MACRO NAND4BX1
    CLASS CORE ;
    FOREIGN NAND4BX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND4BXL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.730 3.000 2.130 3.400 ;
        RECT  2.130 3.000 3.230 3.240 ;
        RECT  3.230 3.000 3.630 3.400 ;
        RECT  3.390 0.920 4.160 1.320 ;
        RECT  3.630 3.000 4.170 3.240 ;
        RECT  4.160 0.920 4.170 1.530 ;
        RECT  4.170 0.920 4.410 3.240 ;
        RECT  4.410 0.920 4.420 1.530 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.440 1.600 1.520 2.000 ;
        RECT  1.520 1.600 1.780 2.090 ;
        RECT  1.780 1.600 1.840 2.000 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.910 2.380 2.500 2.680 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.320 3.240 2.720 ;
        RECT  3.240 2.380 3.760 2.660 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.760 1.720 0.860 2.120 ;
        RECT  0.860 1.720 1.120 2.650 ;
        RECT  1.120 1.720 1.160 2.120 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.040 5.440 ;
        RECT  1.040 4.480 1.440 5.440 ;
        RECT  1.440 4.640 2.420 5.440 ;
        RECT  2.420 4.480 2.820 5.440 ;
        RECT  2.820 4.640 3.940 5.440 ;
        RECT  3.940 4.480 4.340 5.440 ;
        RECT  4.340 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.190 0.400 ;
        RECT  1.190 -0.400 1.590 0.560 ;
        RECT  1.590 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.160 1.600 3.560 2.000 ;
        RECT  3.110 1.600 3.160 1.840 ;
        RECT  2.870 1.080 3.110 1.840 ;
        RECT  0.710 1.080 2.870 1.320 ;
        RECT  0.480 1.040 0.710 1.440 ;
        RECT  0.480 2.930 0.570 3.330 ;
        RECT  0.310 1.040 0.480 3.330 ;
        RECT  0.240 1.120 0.310 3.330 ;
        RECT  0.170 2.930 0.240 3.330 ;
    END
END NAND4BX1

MACRO NAND4XL
    CLASS CORE ;
    FOREIGN NAND4XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.850 3.000 1.250 3.400 ;
        RECT  1.250 3.000 2.350 3.240 ;
        RECT  2.350 3.000 2.750 3.400 ;
        RECT  2.560 0.920 2.960 1.320 ;
        RECT  2.960 1.080 3.500 1.320 ;
        RECT  2.750 3.000 3.510 3.240 ;
        RECT  3.500 1.080 3.510 1.530 ;
        RECT  3.510 1.080 3.750 3.240 ;
        RECT  3.750 1.080 3.760 1.530 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.500 0.460 2.090 ;
        RECT  0.460 1.500 1.000 2.000 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 0.980 2.650 ;
        RECT  0.980 2.390 1.130 2.720 ;
        RECT  1.130 2.320 1.530 2.720 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.850 2.320 2.250 2.720 ;
        RECT  2.250 2.390 2.440 2.650 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.310 1.600 2.710 2.000 ;
        RECT  2.710 1.760 2.840 2.000 ;
        RECT  2.840 1.760 3.100 2.090 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.540 5.440 ;
        RECT  1.540 4.480 1.940 5.440 ;
        RECT  1.940 4.640 3.060 5.440 ;
        RECT  3.060 4.480 3.460 5.440 ;
        RECT  3.460 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.360 0.400 ;
        RECT  0.360 -0.400 0.760 0.560 ;
        RECT  0.760 -0.400 3.960 0.400 ;
        END
    END GND
END NAND4XL

MACRO NAND4X4
    CLASS CORE ;
    FOREIGN NAND4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND4XL ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.990 3.600 1.390 4.000 ;
        RECT  1.390 3.600 2.630 3.840 ;
        RECT  2.630 3.600 3.030 4.000 ;
        RECT  2.660 0.670 4.330 0.910 ;
        RECT  4.330 0.670 4.570 1.100 ;
        RECT  3.030 3.600 7.430 3.840 ;
        RECT  7.430 3.600 7.830 4.000 ;
        RECT  7.830 3.600 8.900 3.840 ;
        RECT  8.900 3.440 9.350 3.840 ;
        RECT  9.350 2.380 9.790 3.840 ;
        RECT  9.790 2.380 9.940 2.660 ;
        RECT  4.570 0.860 9.940 1.100 ;
        RECT  9.940 0.860 10.180 2.660 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.260 0.460 2.090 ;
        RECT  0.460 1.260 0.630 2.010 ;
        RECT  0.630 1.190 0.870 2.010 ;
        RECT  0.870 1.190 3.670 1.430 ;
        RECT  3.670 1.190 3.910 1.620 ;
        RECT  3.910 1.380 4.880 1.620 ;
        RECT  4.880 1.380 5.280 2.010 ;
        RECT  5.280 1.380 9.260 1.620 ;
        RECT  9.260 1.380 9.660 2.010 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.190 2.280 1.350 2.680 ;
        RECT  1.350 2.280 1.590 3.320 ;
        RECT  1.590 2.950 1.780 3.320 ;
        RECT  1.780 3.080 4.430 3.320 ;
        RECT  4.430 2.920 4.830 3.320 ;
        RECT  4.830 2.920 5.630 3.160 ;
        RECT  5.630 2.920 6.270 3.320 ;
        RECT  6.270 2.920 8.510 3.160 ;
        RECT  8.510 2.280 8.750 3.160 ;
        RECT  8.750 2.280 8.910 2.680 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.960 2.260 2.360 2.660 ;
        RECT  2.360 2.390 2.440 2.650 ;
        RECT  2.440 2.410 3.630 2.650 ;
        RECT  3.630 2.290 3.720 2.650 ;
        RECT  3.720 2.290 4.170 2.800 ;
        RECT  4.170 2.290 6.350 2.530 ;
        RECT  6.350 2.040 6.750 2.530 ;
        RECT  6.750 2.290 7.770 2.530 ;
        RECT  7.770 2.120 8.170 2.530 ;
        RECT  8.170 2.200 8.180 2.530 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.790 1.730 3.280 2.100 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 3.820 0.570 5.440 ;
        RECT  0.570 4.640 1.810 5.440 ;
        RECT  1.810 4.480 2.210 5.440 ;
        RECT  2.210 4.640 3.380 5.440 ;
        RECT  3.380 4.300 3.390 5.440 ;
        RECT  3.390 4.180 3.790 5.440 ;
        RECT  3.790 4.300 3.800 5.440 ;
        RECT  3.800 4.640 6.660 5.440 ;
        RECT  6.660 4.300 6.670 5.440 ;
        RECT  6.670 4.180 7.070 5.440 ;
        RECT  7.070 4.300 7.080 5.440 ;
        RECT  7.080 4.640 8.250 5.440 ;
        RECT  8.250 4.480 8.650 5.440 ;
        RECT  8.650 4.640 9.820 5.440 ;
        RECT  9.820 4.320 9.830 5.440 ;
        RECT  9.830 4.120 10.230 5.440 ;
        RECT  10.230 4.320 10.240 5.440 ;
        RECT  10.240 4.640 10.560 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.460 0.400 ;
        RECT  0.460 -0.400 0.860 0.560 ;
        RECT  0.860 -0.400 4.860 0.400 ;
        RECT  4.860 -0.400 5.260 0.560 ;
        RECT  5.260 -0.400 9.260 0.400 ;
        RECT  9.260 -0.400 9.660 0.560 ;
        RECT  9.660 -0.400 10.560 0.400 ;
        END
    END GND
END NAND4X4

MACRO NAND4X2
    CLASS CORE ;
    FOREIGN NAND4X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND4XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.970 0.700 3.510 1.100 ;
        RECT  3.510 0.860 4.730 1.100 ;
        RECT  4.730 0.860 4.820 1.510 ;
        RECT  4.820 0.860 4.970 1.530 ;
        RECT  4.970 1.270 5.080 1.530 ;
        RECT  1.040 3.870 5.490 4.110 ;
        RECT  5.490 3.760 5.530 4.110 ;
        RECT  5.080 1.290 5.530 1.530 ;
        RECT  5.530 1.290 5.770 4.110 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.830 2.240 1.070 3.510 ;
        RECT  1.070 2.390 1.120 2.650 ;
        RECT  1.070 3.200 1.210 3.510 ;
        RECT  1.210 3.270 5.010 3.510 ;
        RECT  5.010 1.810 5.250 3.510 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.550 2.090 ;
        RECT  1.550 1.830 1.780 2.990 ;
        RECT  1.780 1.840 1.790 2.990 ;
        RECT  1.790 2.660 1.870 2.990 ;
        RECT  1.870 2.750 4.480 2.990 ;
        RECT  4.480 2.530 4.720 2.990 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.250 2.200 2.660 2.460 ;
        RECT  2.660 2.220 3.680 2.460 ;
        RECT  3.680 2.180 3.850 2.460 ;
        RECT  3.850 1.850 4.090 2.460 ;
        RECT  4.090 1.850 4.160 2.090 ;
        RECT  4.160 1.830 4.420 2.090 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 1.270 2.190 1.530 ;
        RECT  2.190 1.270 2.440 1.620 ;
        RECT  2.440 1.380 2.930 1.620 ;
        RECT  2.930 1.380 3.170 1.940 ;
        RECT  3.170 1.700 3.360 1.940 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.210 5.440 ;
        RECT  0.210 4.480 0.610 5.440 ;
        RECT  0.610 4.640 1.860 5.440 ;
        RECT  1.860 4.480 2.260 5.440 ;
        RECT  2.260 4.640 3.510 5.440 ;
        RECT  3.510 4.480 3.910 5.440 ;
        RECT  3.910 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.760 0.400 ;
        RECT  0.760 -0.400 0.770 1.040 ;
        RECT  0.770 -0.400 1.170 1.240 ;
        RECT  1.170 -0.400 1.180 1.040 ;
        RECT  1.180 -0.400 5.200 0.400 ;
        RECT  5.200 -0.400 5.600 0.560 ;
        RECT  5.600 -0.400 5.940 0.400 ;
        END
    END GND
END NAND4X2

MACRO NAND4X1
    CLASS CORE ;
    FOREIGN NAND4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND4XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.850 3.000 1.250 3.400 ;
        RECT  1.250 3.000 2.350 3.240 ;
        RECT  2.350 3.000 2.750 3.400 ;
        RECT  2.560 0.920 2.960 1.320 ;
        RECT  2.960 1.080 3.500 1.320 ;
        RECT  2.750 3.000 3.510 3.240 ;
        RECT  3.500 1.080 3.510 1.530 ;
        RECT  3.510 1.080 3.750 3.240 ;
        RECT  3.750 1.270 3.760 1.530 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.470 0.460 2.090 ;
        RECT  0.460 1.470 1.000 2.000 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 0.980 2.650 ;
        RECT  0.980 2.390 1.130 2.720 ;
        RECT  1.130 2.320 1.530 2.720 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.850 2.320 2.250 2.720 ;
        RECT  2.250 2.390 2.440 2.650 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.330 1.600 2.730 2.000 ;
        RECT  2.730 1.760 2.840 2.000 ;
        RECT  2.840 1.760 3.090 2.090 ;
        RECT  3.090 1.830 3.100 2.090 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.540 5.440 ;
        RECT  1.540 4.480 1.940 5.440 ;
        RECT  1.940 4.640 3.060 5.440 ;
        RECT  3.060 4.480 3.460 5.440 ;
        RECT  3.460 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.360 0.400 ;
        RECT  0.360 -0.400 0.760 0.560 ;
        RECT  0.760 -0.400 3.960 0.400 ;
        END
    END GND
END NAND4X1

MACRO NAND3BXL
    CLASS CORE ;
    FOREIGN NAND3BXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.770 2.960 2.170 3.940 ;
        RECT  2.170 2.960 3.190 3.200 ;
        RECT  3.190 2.940 3.360 3.220 ;
        RECT  3.320 0.670 3.410 1.070 ;
        RECT  3.360 2.940 3.520 3.540 ;
        RECT  3.410 0.670 3.520 1.280 ;
        RECT  3.520 0.670 3.760 3.540 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.270 1.540 1.530 ;
        RECT  1.540 1.270 1.780 2.150 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 1.610 2.530 2.120 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.750 2.940 1.260 3.290 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.120 5.440 ;
        RECT  1.120 4.480 2.920 5.440 ;
        RECT  2.920 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.380 0.400 ;
        RECT  1.380 -0.400 1.780 0.560 ;
        RECT  1.780 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.000 2.230 3.240 2.670 ;
        RECT  0.800 2.430 3.000 2.670 ;
        RECT  0.560 0.850 0.800 2.670 ;
        RECT  0.510 3.550 0.650 3.950 ;
        RECT  0.400 0.850 0.560 1.250 ;
        RECT  0.510 2.430 0.560 2.670 ;
        RECT  0.270 2.430 0.510 3.950 ;
        RECT  0.250 3.550 0.270 3.950 ;
    END
END NAND3BXL

MACRO NAND3BX4
    CLASS CORE ;
    FOREIGN NAND3BX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND3BXL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.690 3.500 2.090 4.310 ;
        RECT  2.090 3.500 3.210 3.780 ;
        RECT  3.210 3.500 3.610 4.310 ;
        RECT  3.210 0.730 3.610 1.540 ;
        RECT  3.610 3.500 4.730 3.780 ;
        RECT  4.730 3.500 5.130 4.310 ;
        RECT  5.130 3.500 6.310 3.780 ;
        RECT  3.610 1.300 6.380 1.540 ;
        RECT  6.310 3.010 6.710 3.990 ;
        RECT  6.380 1.260 6.710 1.540 ;
        RECT  6.710 0.730 7.110 1.540 ;
        RECT  6.710 3.490 7.370 3.810 ;
        RECT  7.110 1.300 7.370 1.540 ;
        RECT  7.370 1.300 7.610 3.810 ;
        RECT  7.610 1.820 7.810 3.810 ;
        RECT  7.810 2.640 8.250 3.810 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.390 1.780 2.650 ;
        RECT  1.780 2.150 2.180 2.640 ;
        RECT  2.180 2.400 5.370 2.640 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 2.950 2.190 3.210 ;
        RECT  2.190 2.940 2.440 3.210 ;
        RECT  2.440 2.940 5.790 3.180 ;
        RECT  5.790 2.430 6.030 3.180 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.730 1.820 1.130 2.250 ;
        RECT  1.130 1.820 1.210 2.100 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.920 5.440 ;
        RECT  0.920 4.020 0.930 5.440 ;
        RECT  0.930 3.530 1.330 5.440 ;
        RECT  1.330 4.020 1.340 5.440 ;
        RECT  1.340 4.640 2.440 5.440 ;
        RECT  2.440 4.380 2.450 5.440 ;
        RECT  2.450 4.180 2.850 5.440 ;
        RECT  2.850 4.380 2.860 5.440 ;
        RECT  2.860 4.640 3.960 5.440 ;
        RECT  3.960 4.380 3.970 5.440 ;
        RECT  3.970 4.180 4.370 5.440 ;
        RECT  4.370 4.380 4.380 5.440 ;
        RECT  4.380 4.640 5.480 5.440 ;
        RECT  5.480 4.380 5.490 5.440 ;
        RECT  5.490 4.180 5.890 5.440 ;
        RECT  5.890 4.380 5.900 5.440 ;
        RECT  5.900 4.640 6.990 5.440 ;
        RECT  6.990 4.480 7.390 5.440 ;
        RECT  7.390 4.640 8.580 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.470 0.400 ;
        RECT  1.470 -0.400 1.870 0.560 ;
        RECT  1.870 -0.400 4.970 0.400 ;
        RECT  4.970 -0.400 5.370 0.560 ;
        RECT  5.370 -0.400 8.580 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.930 1.860 6.870 2.100 ;
        RECT  2.690 1.310 2.930 2.100 ;
        RECT  1.060 1.310 2.690 1.550 ;
        RECT  1.050 0.790 1.060 1.550 ;
        RECT  0.650 0.670 1.050 1.550 ;
        RECT  0.640 0.790 0.650 1.550 ;
        RECT  0.450 1.310 0.640 1.550 ;
        RECT  0.450 2.940 0.570 3.920 ;
        RECT  0.210 1.310 0.450 3.920 ;
        RECT  0.170 2.940 0.210 3.920 ;
    END
END NAND3BX4

MACRO NAND3BX2
    CLASS CORE ;
    FOREIGN NAND3BX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND3BXL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.770 0.780 3.170 1.180 ;
        RECT  1.870 3.490 3.500 3.730 ;
        RECT  3.500 3.490 3.760 3.770 ;
        RECT  3.760 3.490 4.830 3.730 ;
        RECT  3.170 0.940 4.830 1.180 ;
        RECT  4.830 0.940 5.070 3.730 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.350 2.240 1.510 2.640 ;
        RECT  1.510 2.240 1.750 3.180 ;
        RECT  1.750 2.940 4.160 3.180 ;
        RECT  4.160 2.940 4.310 3.210 ;
        RECT  4.270 1.520 4.310 1.940 ;
        RECT  4.310 1.520 4.420 3.210 ;
        RECT  4.420 1.520 4.550 3.180 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.070 2.240 2.470 2.640 ;
        RECT  2.470 2.400 2.840 2.640 ;
        RECT  2.840 2.390 2.850 2.650 ;
        RECT  2.850 2.390 3.100 2.660 ;
        RECT  3.100 2.400 3.790 2.660 ;
        RECT  3.790 2.260 4.030 2.660 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.740 1.120 3.210 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.040 5.440 ;
        RECT  1.040 3.920 1.050 5.440 ;
        RECT  1.050 3.720 1.450 5.440 ;
        RECT  1.450 3.920 1.460 5.440 ;
        RECT  1.460 4.640 2.690 5.440 ;
        RECT  2.690 4.480 3.090 5.440 ;
        RECT  3.090 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.040 0.400 ;
        RECT  1.040 -0.400 1.050 1.150 ;
        RECT  1.050 -0.400 1.450 1.350 ;
        RECT  1.450 -0.400 1.460 1.150 ;
        RECT  1.460 -0.400 4.510 0.400 ;
        RECT  4.510 -0.400 4.910 0.560 ;
        RECT  4.910 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.000 1.540 3.400 1.940 ;
        RECT  0.620 1.630 3.000 1.870 ;
        RECT  0.400 1.060 0.620 1.870 ;
        RECT  0.400 3.490 0.620 3.890 ;
        RECT  0.220 1.060 0.400 3.890 ;
        RECT  0.160 1.630 0.220 3.890 ;
    END
END NAND3BX2

MACRO NAND3BX1
    CLASS CORE ;
    FOREIGN NAND3BX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND3BXL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.920 3.180 3.330 3.420 ;
        RECT  3.330 3.100 3.500 3.640 ;
        RECT  3.500 2.950 3.510 3.640 ;
        RECT  3.170 0.750 3.510 0.990 ;
        RECT  3.510 0.750 3.750 3.640 ;
        RECT  3.750 2.950 3.760 3.640 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 1.790 1.780 2.090 ;
        RECT  1.780 1.790 2.150 2.030 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.090 2.380 2.620 2.800 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.780 2.140 1.120 2.660 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.240 5.440 ;
        RECT  1.240 4.480 3.020 5.440 ;
        RECT  3.020 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.430 0.400 ;
        RECT  1.430 -0.400 1.830 0.560 ;
        RECT  1.830 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.990 1.270 3.230 1.940 ;
        RECT  0.950 1.270 2.990 1.510 ;
        RECT  0.550 1.110 0.950 1.510 ;
        RECT  0.500 3.090 0.760 3.490 ;
        RECT  0.500 1.270 0.550 1.510 ;
        RECT  0.260 1.270 0.500 3.490 ;
    END
END NAND3BX1

MACRO NAND3XL
    CLASS CORE ;
    FOREIGN NAND3XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.100 2.960 1.500 3.940 ;
        RECT  1.500 2.960 1.530 3.210 ;
        RECT  1.530 2.970 2.530 3.210 ;
        RECT  2.530 2.970 2.690 3.220 ;
        RECT  2.610 0.670 2.750 1.070 ;
        RECT  2.690 2.970 2.840 3.540 ;
        RECT  2.840 2.950 2.850 3.540 ;
        RECT  2.750 0.670 2.850 1.260 ;
        RECT  2.850 0.670 3.090 3.540 ;
        RECT  3.090 2.950 3.100 3.540 ;
        RECT  3.100 3.110 3.110 3.540 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.220 2.090 ;
        RECT  0.220 1.380 0.460 2.090 ;
        RECT  0.460 1.380 0.550 1.820 ;
        RECT  0.550 1.380 0.880 1.620 ;
        RECT  0.880 1.220 1.120 1.620 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.580 1.870 2.100 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 2.210 2.580 2.660 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.080 5.440 ;
        RECT  1.080 4.480 2.260 5.440 ;
        RECT  2.260 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.870 0.400 ;
        RECT  0.870 -0.400 1.270 0.560 ;
        RECT  1.270 -0.400 3.300 0.400 ;
        END
    END GND
END NAND3XL

MACRO NAND3X4
    CLASS CORE ;
    FOREIGN NAND3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND3XL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.050 3.500 1.450 4.310 ;
        RECT  1.450 3.500 2.570 3.780 ;
        RECT  2.570 3.500 2.970 4.310 ;
        RECT  2.610 0.730 3.010 1.540 ;
        RECT  2.970 3.500 4.090 3.740 ;
        RECT  4.090 3.500 4.490 4.310 ;
        RECT  3.010 1.300 5.610 1.540 ;
        RECT  4.490 3.500 5.670 3.740 ;
        RECT  5.610 1.260 6.050 1.540 ;
        RECT  5.670 3.010 6.070 3.990 ;
        RECT  6.070 3.010 6.280 3.250 ;
        RECT  6.050 0.730 6.450 1.540 ;
        RECT  6.280 2.940 6.710 3.250 ;
        RECT  6.710 1.820 6.760 3.250 ;
        RECT  6.450 1.300 6.760 1.540 ;
        RECT  6.760 1.300 7.000 3.250 ;
        RECT  7.000 1.820 7.150 3.250 ;
        RECT  7.150 2.920 7.210 3.250 ;
        RECT  7.210 2.920 7.610 3.900 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 1.120 2.650 ;
        RECT  1.120 2.150 1.520 2.640 ;
        RECT  1.520 2.400 4.690 2.640 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.950 1.530 3.210 ;
        RECT  1.530 2.940 1.780 3.210 ;
        RECT  1.780 2.940 5.130 3.180 ;
        RECT  5.130 2.430 5.370 3.180 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.550 1.860 2.840 2.100 ;
        RECT  2.840 1.830 3.100 2.100 ;
        RECT  3.100 1.860 6.210 2.100 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.020 0.170 5.440 ;
        RECT  0.170 3.820 0.570 5.440 ;
        RECT  0.570 4.020 0.580 5.440 ;
        RECT  0.580 4.640 1.800 5.440 ;
        RECT  1.800 4.380 1.810 5.440 ;
        RECT  1.810 4.180 2.210 5.440 ;
        RECT  2.210 4.380 2.220 5.440 ;
        RECT  2.220 4.640 3.320 5.440 ;
        RECT  3.320 4.180 3.730 5.440 ;
        RECT  3.730 4.380 3.740 5.440 ;
        RECT  3.740 4.640 4.840 5.440 ;
        RECT  4.840 4.380 4.850 5.440 ;
        RECT  4.850 4.180 5.250 5.440 ;
        RECT  5.250 4.380 5.260 5.440 ;
        RECT  5.260 4.640 6.340 5.440 ;
        RECT  6.340 4.480 6.740 5.440 ;
        RECT  6.740 4.640 7.920 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.860 0.400 ;
        RECT  0.860 -0.400 0.870 1.020 ;
        RECT  0.870 -0.400 1.270 1.220 ;
        RECT  1.270 -0.400 1.280 1.020 ;
        RECT  1.280 -0.400 4.300 0.400 ;
        RECT  4.300 -0.400 4.310 0.810 ;
        RECT  4.310 -0.400 4.710 1.010 ;
        RECT  4.710 -0.400 4.720 0.810 ;
        RECT  4.720 -0.400 7.920 0.400 ;
        END
    END GND
END NAND3X4

MACRO NAND3X2
    CLASS CORE ;
    FOREIGN NAND3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND3XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.820 1.130 1.060 3.400 ;
        RECT  1.060 1.130 1.120 1.530 ;
        RECT  1.060 3.000 1.330 3.400 ;
        RECT  1.120 1.130 1.770 1.450 ;
        RECT  1.770 1.040 2.070 1.450 ;
        RECT  2.070 1.050 2.310 1.450 ;
        RECT  1.330 3.080 2.570 3.320 ;
        RECT  2.570 3.000 2.970 3.400 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.210 2.650 ;
        RECT  0.210 2.310 0.300 2.650 ;
        RECT  0.300 2.230 0.540 3.920 ;
        RECT  0.540 3.680 3.490 3.920 ;
        RECT  3.490 1.800 3.730 3.920 ;
        RECT  3.730 1.800 3.890 2.530 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.340 2.240 1.580 2.720 ;
        RECT  1.580 2.480 2.840 2.720 ;
        RECT  2.840 2.390 2.850 2.720 ;
        RECT  2.850 2.240 3.090 2.720 ;
        RECT  3.090 2.390 3.100 2.650 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.010 1.800 2.090 2.200 ;
        RECT  2.090 1.790 2.440 2.210 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.320 0.170 5.440 ;
        RECT  0.170 4.200 0.570 5.440 ;
        RECT  0.570 4.320 0.580 5.440 ;
        RECT  0.580 4.640 1.750 5.440 ;
        RECT  1.750 4.480 2.150 5.440 ;
        RECT  2.150 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 3.590 0.400 ;
        RECT  3.590 -0.400 3.600 1.070 ;
        RECT  3.600 -0.400 4.000 1.270 ;
        RECT  4.000 -0.400 4.010 1.070 ;
        RECT  4.010 -0.400 4.620 0.400 ;
        END
    END GND
END NAND3X2

MACRO NAND3X1
    CLASS CORE ;
    FOREIGN NAND3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND3XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.740 3.100 1.140 3.500 ;
        RECT  1.140 3.180 2.090 3.420 ;
        RECT  2.090 3.180 2.120 3.520 ;
        RECT  2.120 3.090 2.240 3.520 ;
        RECT  2.240 0.860 2.480 3.740 ;
        RECT  2.480 2.950 3.100 3.740 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.210 2.090 ;
        RECT  0.210 1.500 0.560 2.090 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.830 2.380 1.300 2.780 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.270 1.720 1.530 ;
        RECT  1.720 1.270 1.780 2.410 ;
        RECT  1.780 1.280 1.960 2.410 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 1.700 5.440 ;
        RECT  1.700 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 3.300 0.400 ;
        END
    END GND
END NAND3X1

MACRO NAND2BXL
    CLASS CORE ;
    FOREIGN NAND2BXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 1.270 2.210 1.530 ;
        RECT  1.810 3.500 2.650 3.740 ;
        RECT  2.210 1.120 2.650 1.540 ;
        RECT  2.650 1.120 2.890 3.740 ;
        RECT  2.890 1.120 2.900 1.540 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 2.530 1.520 2.940 ;
        RECT  1.520 2.530 1.780 3.210 ;
        RECT  1.780 2.530 1.870 2.940 ;
        RECT  1.870 2.530 1.880 2.930 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.760 2.390 1.120 3.000 ;
        RECT  1.120 2.600 1.160 3.000 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.040 5.440 ;
        RECT  1.040 4.480 1.440 5.440 ;
        RECT  1.440 4.640 2.630 5.440 ;
        RECT  2.630 4.480 3.030 5.440 ;
        RECT  3.030 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.060 0.400 ;
        RECT  1.060 -0.400 1.070 1.290 ;
        RECT  1.070 -0.400 1.470 1.490 ;
        RECT  1.470 -0.400 1.480 1.290 ;
        RECT  1.480 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.130 1.810 2.370 2.210 ;
        RECT  0.590 1.810 2.130 2.050 ;
        RECT  0.480 1.330 0.590 2.050 ;
        RECT  0.480 3.240 0.590 3.640 ;
        RECT  0.240 1.330 0.480 3.640 ;
        RECT  0.190 1.330 0.240 1.730 ;
        RECT  0.190 3.240 0.240 3.640 ;
    END
END NAND2BXL

MACRO NAND2BX4
    CLASS CORE ;
    FOREIGN NAND2BX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND2BXL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.980 2.940 2.380 4.000 ;
        RECT  2.270 1.020 2.670 1.420 ;
        RECT  2.380 2.940 3.410 3.250 ;
        RECT  3.410 2.940 3.850 4.340 ;
        RECT  3.850 2.940 3.900 4.000 ;
        RECT  2.670 1.180 4.710 1.420 ;
        RECT  3.900 2.940 5.060 3.250 ;
        RECT  4.710 1.070 5.060 1.470 ;
        RECT  5.060 1.070 5.110 3.250 ;
        RECT  5.110 1.150 5.300 3.250 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.410 1.690 1.650 2.090 ;
        RECT  1.650 1.720 1.780 2.090 ;
        RECT  1.780 1.720 3.690 1.960 ;
        RECT  3.690 1.700 4.090 2.100 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.160 1.830 0.600 2.470 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.210 5.440 ;
        RECT  1.210 4.370 1.220 5.440 ;
        RECT  1.220 4.170 1.620 5.440 ;
        RECT  1.620 4.370 1.630 5.440 ;
        RECT  1.630 4.640 2.730 5.440 ;
        RECT  2.730 4.090 2.740 5.440 ;
        RECT  2.740 3.600 3.140 5.440 ;
        RECT  3.140 4.090 3.150 5.440 ;
        RECT  3.150 4.640 4.310 5.440 ;
        RECT  4.310 4.020 4.320 5.440 ;
        RECT  4.320 3.820 4.720 5.440 ;
        RECT  4.720 4.020 4.730 5.440 ;
        RECT  4.730 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.020 0.400 ;
        RECT  1.020 -0.400 1.030 0.660 ;
        RECT  1.030 -0.400 1.430 0.780 ;
        RECT  1.430 -0.400 1.440 0.660 ;
        RECT  1.440 -0.400 3.480 0.400 ;
        RECT  3.480 -0.400 3.490 0.670 ;
        RECT  3.490 -0.400 3.890 0.790 ;
        RECT  3.890 -0.400 3.900 0.670 ;
        RECT  3.900 -0.400 5.940 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.540 2.070 4.780 2.640 ;
        RECT  2.890 2.400 4.540 2.640 ;
        RECT  2.490 2.240 2.890 2.640 ;
        RECT  1.130 2.400 2.490 2.640 ;
        RECT  0.890 1.250 1.130 3.730 ;
        RECT  0.870 1.250 0.890 2.640 ;
        RECT  0.760 3.490 0.890 3.730 ;
        RECT  0.670 1.250 0.870 1.490 ;
        RECT  0.360 3.490 0.760 3.890 ;
        RECT  0.270 1.090 0.670 1.490 ;
    END
END NAND2BX4

MACRO NAND2BX2
    CLASS CORE ;
    FOREIGN NAND2BX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND2BXL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.570 3.000 2.840 3.240 ;
        RECT  2.840 2.950 3.100 3.240 ;
        RECT  3.100 3.000 3.710 3.240 ;
        RECT  2.270 1.270 3.710 1.510 ;
        RECT  3.710 1.270 3.950 3.240 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.350 2.400 1.520 2.640 ;
        RECT  1.520 2.390 1.780 2.650 ;
        RECT  1.780 2.400 3.190 2.640 ;
        RECT  3.190 2.240 3.430 2.640 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.860 0.460 2.650 ;
        RECT  0.460 1.860 0.490 2.380 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.550 5.440 ;
        RECT  1.550 4.480 1.890 5.440 ;
        RECT  1.890 4.450 3.080 5.440 ;
        RECT  3.080 4.480 3.410 5.440 ;
        RECT  3.410 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        RECT  0.990 -0.400 1.390 0.560 ;
        RECT  1.390 -0.400 3.550 0.400 ;
        RECT  3.550 -0.400 3.950 0.560 ;
        RECT  3.950 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.060 1.870 2.670 2.110 ;
        RECT  0.820 1.300 1.060 3.740 ;
        RECT  0.570 1.300 0.820 1.550 ;
        RECT  0.170 3.500 0.820 3.740 ;
        RECT  0.170 1.140 0.570 1.550 ;
    END
END NAND2BX2

MACRO NAND2BX1
    CLASS CORE ;
    FOREIGN NAND2BX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND2BXL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.810 3.500 2.800 3.740 ;
        RECT  2.180 1.170 2.800 1.590 ;
        RECT  2.800 1.170 3.040 3.740 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 2.530 1.520 2.940 ;
        RECT  1.520 2.530 1.780 3.210 ;
        RECT  1.780 2.530 1.870 2.940 ;
        RECT  1.870 2.530 1.880 2.930 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.760 2.380 1.210 2.790 ;
        END
    END AN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.040 5.440 ;
        RECT  1.040 4.480 1.440 5.440 ;
        RECT  1.440 4.640 2.630 5.440 ;
        RECT  2.630 4.480 3.030 5.440 ;
        RECT  3.030 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.060 0.400 ;
        RECT  1.060 -0.400 1.070 1.290 ;
        RECT  1.070 -0.400 1.470 1.490 ;
        RECT  1.470 -0.400 1.480 1.290 ;
        RECT  1.480 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.280 1.860 2.520 2.320 ;
        RECT  0.590 1.860 2.280 2.100 ;
        RECT  0.480 1.350 0.590 2.100 ;
        RECT  0.480 3.110 0.590 3.510 ;
        RECT  0.240 1.350 0.480 3.510 ;
        RECT  0.190 1.350 0.240 1.750 ;
        RECT  0.190 3.110 0.240 3.510 ;
    END
END NAND2BX1

MACRO NAND2XL
    CLASS CORE ;
    FOREIGN NAND2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.840 3.120 0.850 3.540 ;
        RECT  0.850 3.090 1.520 3.540 ;
        RECT  1.520 2.950 1.570 3.540 ;
        RECT  1.370 1.150 1.570 1.550 ;
        RECT  1.570 1.150 1.810 3.540 ;
        RECT  1.810 3.120 1.820 3.540 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.180 1.960 0.510 2.650 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 1.050 2.090 ;
        RECT  1.050 1.830 1.120 2.670 ;
        RECT  1.120 1.840 1.290 2.670 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 1.980 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.980 0.400 ;
        END
    END GND
END NAND2XL

MACRO NAND2X4
    CLASS CORE ;
    FOREIGN NAND2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND2XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.770 2.940 1.210 4.340 ;
        RECT  1.210 2.940 1.330 3.940 ;
        RECT  1.450 0.770 1.850 1.170 ;
        RECT  1.330 2.940 2.450 3.220 ;
        RECT  2.450 2.940 2.850 3.940 ;
        RECT  2.850 2.940 2.980 3.190 ;
        RECT  1.850 0.860 3.630 1.100 ;
        RECT  3.630 0.850 4.010 1.100 ;
        RECT  2.980 2.950 4.090 3.190 ;
        RECT  4.010 0.850 4.090 1.400 ;
        RECT  4.090 0.850 4.330 3.190 ;
        RECT  4.330 0.850 4.410 1.400 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.060 0.890 2.660 ;
        RECT  0.890 2.380 2.680 2.660 ;
        RECT  2.680 2.250 2.740 2.660 ;
        RECT  2.740 2.240 3.090 2.660 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.510 1.730 1.910 2.110 ;
        RECT  1.910 1.730 3.570 1.970 ;
        RECT  3.570 1.730 3.810 2.470 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.250 5.440 ;
        RECT  0.250 3.540 0.490 5.440 ;
        RECT  0.490 4.640 1.680 5.440 ;
        RECT  1.680 4.030 1.690 5.440 ;
        RECT  1.690 3.540 2.090 5.440 ;
        RECT  2.090 4.030 2.100 5.440 ;
        RECT  2.100 4.640 3.260 5.440 ;
        RECT  3.260 4.020 3.270 5.440 ;
        RECT  3.270 3.820 3.670 5.440 ;
        RECT  3.670 4.020 3.680 5.440 ;
        RECT  3.680 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 2.730 0.400 ;
        RECT  2.730 -0.400 3.130 0.560 ;
        RECT  3.130 -0.400 5.280 0.400 ;
        END
    END GND
END NAND2X4

MACRO NAND2X2
    CLASS CORE ;
    FOREIGN NAND2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND2XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.750 2.940 1.150 3.350 ;
        RECT  1.450 1.050 1.850 1.450 ;
        RECT  1.150 2.940 2.130 3.220 ;
        RECT  1.850 1.210 2.210 1.450 ;
        RECT  2.210 1.210 2.450 1.870 ;
        RECT  2.130 2.940 2.530 3.350 ;
        RECT  2.530 2.940 2.890 3.220 ;
        RECT  2.450 1.630 2.890 1.870 ;
        RECT  2.890 1.630 3.130 3.220 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.480 2.250 0.770 2.650 ;
        RECT  0.770 2.250 0.880 2.660 ;
        RECT  0.880 2.390 1.540 2.660 ;
        RECT  1.540 2.390 2.370 2.630 ;
        RECT  2.370 2.220 2.610 2.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.390 1.740 1.870 2.120 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.470 5.440 ;
        RECT  1.470 4.480 1.870 5.440 ;
        RECT  1.870 4.640 2.730 5.440 ;
        RECT  2.730 4.480 3.130 5.440 ;
        RECT  3.130 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.220 0.400 ;
        RECT  0.220 -0.400 0.230 1.210 ;
        RECT  0.230 -0.400 0.630 1.410 ;
        RECT  0.630 -0.400 0.640 1.210 ;
        RECT  0.640 -0.400 2.720 0.400 ;
        RECT  2.720 -0.400 2.730 1.150 ;
        RECT  2.730 -0.400 3.130 1.350 ;
        RECT  3.130 -0.400 3.140 1.150 ;
        RECT  3.140 -0.400 3.300 0.400 ;
        END
    END GND
END NAND2X2

MACRO NAND2X1
    CLASS CORE ;
    FOREIGN NAND2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ NAND2XL ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.770 3.060 1.170 3.460 ;
        RECT  1.230 1.400 1.430 1.800 ;
        RECT  1.170 3.060 1.570 3.300 ;
        RECT  1.430 1.400 1.570 2.090 ;
        RECT  1.570 1.400 1.810 3.300 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.190 1.820 0.490 2.490 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.360 1.120 2.780 ;
        RECT  1.120 2.370 1.290 2.770 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.460 0.570 5.440 ;
        RECT  0.570 4.640 1.410 5.440 ;
        RECT  1.410 4.480 1.810 5.440 ;
        RECT  1.810 4.640 1.980 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.980 0.400 ;
        END
    END GND
END NAND2X1

MACRO MXI4XL
    CLASS CORE ;
    FOREIGN MXI4XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.520 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.130 3.930 13.530 4.370 ;
        RECT  13.530 3.930 13.970 4.170 ;
        RECT  13.710 1.390 13.970 1.790 ;
        RECT  13.970 1.390 14.110 4.170 ;
        RECT  14.110 1.550 14.210 4.170 ;
        RECT  14.210 2.390 14.320 2.650 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  12.620 2.250 13.090 2.660 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.110 2.210 4.530 2.660 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.400 1.270 5.820 2.020 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.290 1.610 8.690 2.070 ;
        RECT  8.690 1.830 8.780 2.070 ;
        RECT  8.780 1.830 9.040 2.090 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.280 1.660 3.500 2.080 ;
        RECT  3.500 1.660 3.680 2.090 ;
        RECT  3.680 1.830 3.760 2.090 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.460 2.470 ;
        RECT  0.460 1.840 0.800 2.470 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 3.610 5.440 ;
        RECT  3.610 4.110 3.620 5.440 ;
        RECT  3.620 3.990 4.020 5.440 ;
        RECT  4.020 4.110 4.030 5.440 ;
        RECT  4.030 4.640 5.230 5.440 ;
        RECT  5.230 4.110 5.240 5.440 ;
        RECT  5.240 3.990 5.640 5.440 ;
        RECT  5.640 4.110 5.650 5.440 ;
        RECT  5.650 4.640 8.500 5.440 ;
        RECT  8.500 4.480 8.900 5.440 ;
        RECT  8.900 4.640 12.040 5.440 ;
        RECT  12.040 3.650 12.050 5.440 ;
        RECT  12.050 3.450 12.450 5.440 ;
        RECT  12.450 3.650 12.460 5.440 ;
        RECT  12.460 4.640 13.950 5.440 ;
        RECT  13.950 4.480 14.350 5.440 ;
        RECT  14.350 4.640 14.520 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 3.450 0.400 ;
        RECT  3.450 -0.400 3.460 1.180 ;
        RECT  3.460 -0.400 3.860 1.380 ;
        RECT  3.860 -0.400 3.870 1.180 ;
        RECT  3.870 -0.400 5.260 0.400 ;
        RECT  5.260 -0.400 5.270 0.860 ;
        RECT  5.270 -0.400 5.670 0.980 ;
        RECT  5.670 -0.400 5.680 0.860 ;
        RECT  5.680 -0.400 8.500 0.400 ;
        RECT  8.500 -0.400 8.900 0.560 ;
        RECT  8.900 -0.400 11.960 0.400 ;
        RECT  11.960 -0.400 11.970 0.750 ;
        RECT  11.970 -0.400 12.370 0.870 ;
        RECT  12.370 -0.400 12.380 0.750 ;
        RECT  12.380 -0.400 13.710 0.400 ;
        RECT  13.710 -0.400 14.110 0.560 ;
        RECT  14.110 -0.400 14.520 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  13.240 0.670 13.400 0.910 ;
        RECT  13.180 3.190 13.340 3.590 ;
        RECT  12.380 1.670 13.260 1.910 ;
        RECT  13.000 0.670 13.240 1.390 ;
        RECT  12.940 2.930 13.180 3.590 ;
        RECT  11.690 1.150 13.000 1.390 ;
        RECT  12.380 2.930 12.940 3.170 ;
        RECT  12.140 1.670 12.380 3.170 ;
        RECT  11.770 1.670 12.140 1.910 ;
        RECT  11.770 2.650 11.860 3.050 ;
        RECT  11.530 1.670 11.770 2.150 ;
        RECT  11.530 2.650 11.770 4.180 ;
        RECT  11.450 0.670 11.690 1.390 ;
        RECT  11.430 1.910 11.530 2.150 ;
        RECT  6.590 3.940 11.530 4.180 ;
        RECT  10.390 0.670 11.450 0.910 ;
        RECT  11.190 1.910 11.430 2.330 ;
        RECT  10.910 3.030 11.250 3.430 ;
        RECT  10.930 1.190 11.170 1.590 ;
        RECT  10.910 1.350 10.930 1.590 ;
        RECT  10.670 1.350 10.910 3.430 ;
        RECT  10.150 0.670 10.390 3.570 ;
        RECT  9.640 1.140 9.710 1.540 ;
        RECT  9.640 3.030 9.710 3.430 ;
        RECT  9.400 1.140 9.640 3.430 ;
        RECT  9.310 1.140 9.400 1.540 ;
        RECT  9.310 3.030 9.400 3.430 ;
        RECT  8.530 2.410 9.120 2.650 ;
        RECT  8.290 2.410 8.530 3.570 ;
        RECT  7.490 3.330 8.290 3.570 ;
        RECT  7.770 0.990 8.010 3.050 ;
        RECT  7.250 1.020 7.490 3.570 ;
        RECT  6.930 1.020 7.250 1.260 ;
        RECT  6.870 3.330 7.250 3.570 ;
        RECT  6.730 1.610 6.970 3.050 ;
        RECT  6.570 1.610 6.730 1.850 ;
        RECT  6.510 2.810 6.730 3.050 ;
        RECT  6.350 3.470 6.590 4.180 ;
        RECT  6.330 0.990 6.570 1.850 ;
        RECT  6.110 2.810 6.510 3.190 ;
        RECT  6.210 2.130 6.450 2.530 ;
        RECT  2.200 3.470 6.350 3.710 ;
        RECT  6.170 0.990 6.330 1.390 ;
        RECT  5.040 2.290 6.210 2.530 ;
        RECT  4.800 1.410 5.040 3.170 ;
        RECT  4.740 1.410 4.800 1.650 ;
        RECT  3.590 2.930 4.800 3.170 ;
        RECT  4.340 1.250 4.740 1.650 ;
        RECT  3.350 2.370 3.590 3.170 ;
        RECT  2.880 2.370 3.350 2.610 ;
        RECT  2.360 2.890 3.040 3.130 ;
        RECT  2.820 1.060 2.980 1.460 ;
        RECT  2.640 2.210 2.880 2.610 ;
        RECT  2.580 1.060 2.820 1.850 ;
        RECT  2.360 1.610 2.580 1.850 ;
        RECT  2.120 1.610 2.360 3.130 ;
        RECT  1.840 1.090 2.200 1.330 ;
        RECT  1.880 3.410 2.200 3.710 ;
        RECT  1.840 3.410 1.880 3.650 ;
        RECT  1.600 1.090 1.840 3.650 ;
        RECT  1.080 1.040 1.320 3.460 ;
    END
END MXI4XL

MACRO MXI4X4
    CLASS CORE ;
    FOREIGN MXI4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MXI4XL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.170 2.840 15.290 3.820 ;
        RECT  15.170 0.670 15.290 1.650 ;
        RECT  15.290 0.670 15.570 3.820 ;
        RECT  15.570 0.680 15.580 3.220 ;
        RECT  15.580 1.820 15.730 3.220 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  12.080 1.830 12.090 2.090 ;
        RECT  12.090 1.830 12.550 2.230 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.980 1.840 4.160 2.280 ;
        RECT  4.160 1.830 4.380 2.280 ;
        RECT  4.380 1.830 4.420 2.090 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.820 2.160 5.170 2.670 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.310 1.960 8.450 2.360 ;
        RECT  8.450 1.290 8.690 2.360 ;
        RECT  8.690 1.290 8.780 1.530 ;
        RECT  8.780 1.270 9.040 1.530 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.260 2.040 3.420 2.280 ;
        RECT  3.420 1.280 3.500 2.280 ;
        RECT  3.500 1.270 3.660 2.280 ;
        RECT  3.660 1.270 3.760 1.530 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.020 0.790 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.190 5.440 ;
        RECT  0.190 3.690 0.200 5.440 ;
        RECT  0.200 3.490 0.600 5.440 ;
        RECT  0.600 3.690 0.610 5.440 ;
        RECT  0.610 4.640 3.550 5.440 ;
        RECT  3.550 4.240 3.560 5.440 ;
        RECT  3.560 4.120 3.960 5.440 ;
        RECT  3.960 4.240 3.970 5.440 ;
        RECT  3.970 4.640 5.120 5.440 ;
        RECT  5.120 4.240 5.130 5.440 ;
        RECT  5.130 4.120 5.530 5.440 ;
        RECT  5.530 4.240 5.540 5.440 ;
        RECT  5.540 4.640 8.650 5.440 ;
        RECT  8.650 4.480 9.050 5.440 ;
        RECT  9.050 4.640 11.850 5.440 ;
        RECT  11.850 4.480 13.190 5.440 ;
        RECT  13.190 4.640 14.350 5.440 ;
        RECT  14.350 4.480 14.750 5.440 ;
        RECT  14.750 4.640 15.920 5.440 ;
        RECT  15.920 4.080 15.930 5.440 ;
        RECT  15.930 3.590 16.330 5.440 ;
        RECT  16.330 4.080 16.340 5.440 ;
        RECT  16.340 4.640 16.500 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.190 0.400 ;
        RECT  0.190 -0.400 0.200 0.980 ;
        RECT  0.200 -0.400 0.600 1.180 ;
        RECT  0.600 -0.400 0.610 0.980 ;
        RECT  0.610 -0.400 3.550 0.400 ;
        RECT  3.550 -0.400 3.560 0.870 ;
        RECT  3.560 -0.400 3.960 0.990 ;
        RECT  3.960 -0.400 3.970 0.870 ;
        RECT  3.970 -0.400 5.120 0.400 ;
        RECT  5.120 -0.400 5.130 0.860 ;
        RECT  5.130 -0.400 5.530 0.980 ;
        RECT  5.530 -0.400 5.540 0.860 ;
        RECT  5.540 -0.400 8.520 0.400 ;
        RECT  8.520 -0.400 8.530 0.790 ;
        RECT  8.530 -0.400 8.930 0.990 ;
        RECT  8.930 -0.400 8.940 0.790 ;
        RECT  8.940 -0.400 12.770 0.400 ;
        RECT  12.770 -0.400 13.170 0.560 ;
        RECT  13.170 -0.400 14.350 0.400 ;
        RECT  14.350 -0.400 14.750 0.560 ;
        RECT  14.750 -0.400 15.920 0.400 ;
        RECT  15.920 -0.400 15.930 1.070 ;
        RECT  15.930 -0.400 16.330 1.560 ;
        RECT  16.330 -0.400 16.340 1.070 ;
        RECT  16.340 -0.400 16.500 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.860 1.930 15.020 2.330 ;
        RECT  14.620 0.860 14.860 2.330 ;
        RECT  12.490 0.860 14.620 1.100 ;
        RECT  14.210 2.610 14.450 4.180 ;
        RECT  13.920 2.610 14.210 2.850 ;
        RECT  6.210 3.940 14.210 4.180 ;
        RECT  13.230 1.380 13.990 1.620 ;
        RECT  13.230 3.190 13.930 3.660 ;
        RECT  13.680 2.110 13.920 2.850 ;
        RECT  13.520 2.110 13.680 2.510 ;
        RECT  12.990 1.380 13.230 3.660 ;
        RECT  11.410 3.420 12.990 3.660 ;
        RECT  12.250 0.680 12.490 1.100 ;
        RECT  11.990 2.670 12.390 3.140 ;
        RECT  10.470 0.680 12.250 0.920 ;
        RECT  11.720 2.670 11.990 2.910 ;
        RECT  11.720 1.320 11.970 1.560 ;
        RECT  11.480 1.320 11.720 2.910 ;
        RECT  11.430 1.820 11.480 2.220 ;
        RECT  11.070 3.260 11.410 3.660 ;
        RECT  11.070 1.200 11.150 1.600 ;
        RECT  10.830 1.200 11.070 3.660 ;
        RECT  10.470 3.030 10.550 3.430 ;
        RECT  10.230 0.680 10.470 3.430 ;
        RECT  10.070 1.050 10.230 1.450 ;
        RECT  9.550 0.750 9.790 3.430 ;
        RECT  9.310 0.750 9.550 0.990 ;
        RECT  9.030 2.030 9.270 3.660 ;
        RECT  7.510 3.420 9.030 3.660 ;
        RECT  7.790 1.140 8.030 3.140 ;
        RECT  7.270 0.950 7.510 3.660 ;
        RECT  6.950 0.950 7.270 1.350 ;
        RECT  6.710 3.420 7.270 3.660 ;
        RECT  6.750 1.630 6.990 3.070 ;
        RECT  6.590 1.630 6.750 1.870 ;
        RECT  6.270 2.830 6.750 3.070 ;
        RECT  6.350 1.030 6.590 1.870 ;
        RECT  5.680 2.150 6.470 2.550 ;
        RECT  6.190 1.030 6.350 1.430 ;
        RECT  6.030 2.830 6.270 3.240 ;
        RECT  5.970 3.600 6.210 4.180 ;
        RECT  1.820 3.600 5.970 3.840 ;
        RECT  5.440 1.260 5.680 3.180 ;
        RECT  4.780 1.260 5.440 1.500 ;
        RECT  4.440 2.940 5.440 3.180 ;
        RECT  4.380 1.060 4.780 1.500 ;
        RECT  4.200 2.560 4.440 3.180 ;
        RECT  2.860 2.560 4.200 2.800 ;
        RECT  2.890 1.060 3.050 1.460 ;
        RECT  2.340 3.080 2.980 3.320 ;
        RECT  2.650 1.060 2.890 1.850 ;
        RECT  2.620 2.180 2.860 2.800 ;
        RECT  2.340 1.610 2.650 1.850 ;
        RECT  2.100 1.610 2.340 3.320 ;
        RECT  1.820 0.930 2.180 1.330 ;
        RECT  1.580 0.930 1.820 3.840 ;
        RECT  1.060 0.990 1.300 3.460 ;
    END
END MXI4X4

MACRO MXI4X2
    CLASS CORE ;
    FOREIGN MXI4X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MXI4XL ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.720 2.950 14.830 3.210 ;
        RECT  14.830 2.940 15.240 3.210 ;
        RECT  15.240 2.810 15.380 3.210 ;
        RECT  15.250 0.860 15.380 1.400 ;
        RECT  15.380 0.860 15.620 3.210 ;
        RECT  15.620 2.510 15.640 3.210 ;
        RECT  15.620 0.860 15.650 1.400 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  11.990 1.830 12.550 2.230 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.980 1.840 4.160 2.370 ;
        RECT  4.160 1.830 4.380 2.370 ;
        RECT  4.380 1.830 4.420 2.090 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.420 1.270 5.430 1.850 ;
        RECT  5.430 1.270 5.830 2.040 ;
        RECT  5.830 1.270 5.840 1.850 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.310 1.960 8.450 2.360 ;
        RECT  8.450 1.290 8.690 2.360 ;
        RECT  8.690 1.290 8.780 1.530 ;
        RECT  8.780 1.270 9.040 1.530 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.260 1.860 3.420 2.100 ;
        RECT  3.420 1.280 3.500 2.100 ;
        RECT  3.500 1.270 3.660 2.100 ;
        RECT  3.660 1.270 3.760 1.530 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.000 0.790 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.190 5.440 ;
        RECT  0.190 3.690 0.200 5.440 ;
        RECT  0.200 3.490 0.600 5.440 ;
        RECT  0.600 3.690 0.610 5.440 ;
        RECT  0.610 4.640 3.550 5.440 ;
        RECT  3.550 4.060 3.560 5.440 ;
        RECT  3.560 3.940 3.960 5.440 ;
        RECT  3.960 4.060 3.970 5.440 ;
        RECT  3.970 4.640 5.120 5.440 ;
        RECT  5.120 4.060 5.130 5.440 ;
        RECT  5.130 3.940 5.530 5.440 ;
        RECT  5.530 4.060 5.540 5.440 ;
        RECT  5.540 4.640 8.650 5.440 ;
        RECT  8.650 4.480 9.050 5.440 ;
        RECT  9.050 4.640 12.490 5.440 ;
        RECT  12.490 4.480 12.890 5.440 ;
        RECT  12.890 4.640 14.400 5.440 ;
        RECT  14.400 4.480 14.800 5.440 ;
        RECT  14.800 4.640 15.840 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.190 0.400 ;
        RECT  0.190 -0.400 0.200 0.980 ;
        RECT  0.200 -0.400 0.600 1.180 ;
        RECT  0.600 -0.400 0.610 0.980 ;
        RECT  0.610 -0.400 3.550 0.400 ;
        RECT  3.550 -0.400 3.560 0.870 ;
        RECT  3.560 -0.400 3.960 0.990 ;
        RECT  3.960 -0.400 3.970 0.870 ;
        RECT  3.970 -0.400 5.360 0.400 ;
        RECT  5.360 -0.400 5.370 0.860 ;
        RECT  5.370 -0.400 5.770 0.980 ;
        RECT  5.770 -0.400 5.780 0.860 ;
        RECT  5.780 -0.400 8.530 0.400 ;
        RECT  8.530 -0.400 8.930 0.980 ;
        RECT  8.930 -0.400 12.770 0.400 ;
        RECT  12.770 -0.400 13.170 0.560 ;
        RECT  13.170 -0.400 14.430 0.400 ;
        RECT  14.430 -0.400 14.830 0.560 ;
        RECT  14.830 -0.400 15.840 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.770 1.800 15.140 2.200 ;
        RECT  14.740 0.860 14.770 2.200 ;
        RECT  14.530 0.860 14.740 2.120 ;
        RECT  12.490 0.860 14.530 1.100 ;
        RECT  14.010 2.280 14.250 4.180 ;
        RECT  13.240 1.380 14.050 1.620 ;
        RECT  13.920 2.280 14.010 2.520 ;
        RECT  6.210 3.940 14.010 4.180 ;
        RECT  13.520 2.120 13.920 2.520 ;
        RECT  13.240 3.190 13.730 3.590 ;
        RECT  13.000 1.380 13.240 3.590 ;
        RECT  11.410 3.350 13.000 3.590 ;
        RECT  12.250 0.680 12.490 1.100 ;
        RECT  11.950 2.670 12.350 3.070 ;
        RECT  10.470 0.680 12.250 0.920 ;
        RECT  11.720 1.300 11.970 1.540 ;
        RECT  11.720 2.670 11.950 2.910 ;
        RECT  11.480 1.300 11.720 2.910 ;
        RECT  11.350 1.910 11.480 2.310 ;
        RECT  11.070 3.190 11.410 3.590 ;
        RECT  11.070 1.200 11.150 1.600 ;
        RECT  10.830 1.200 11.070 3.590 ;
        RECT  10.390 3.030 10.550 3.430 ;
        RECT  10.390 0.680 10.470 1.330 ;
        RECT  10.230 0.680 10.390 3.430 ;
        RECT  10.150 0.930 10.230 3.430 ;
        RECT  10.070 0.930 10.150 1.330 ;
        RECT  9.550 0.750 9.790 3.430 ;
        RECT  9.310 0.750 9.550 0.990 ;
        RECT  9.030 2.220 9.270 3.600 ;
        RECT  7.510 3.360 9.030 3.600 ;
        RECT  7.790 1.010 8.030 3.070 ;
        RECT  7.270 0.950 7.510 3.600 ;
        RECT  6.950 0.950 7.270 1.350 ;
        RECT  6.710 3.360 7.270 3.600 ;
        RECT  6.750 1.630 6.990 3.080 ;
        RECT  6.590 1.630 6.750 1.870 ;
        RECT  6.350 2.840 6.750 3.080 ;
        RECT  6.350 1.030 6.590 1.870 ;
        RECT  6.230 2.150 6.470 2.560 ;
        RECT  6.190 1.030 6.350 1.430 ;
        RECT  5.950 2.840 6.350 3.130 ;
        RECT  5.020 2.320 6.230 2.560 ;
        RECT  5.970 3.420 6.210 4.180 ;
        RECT  1.820 3.420 5.970 3.660 ;
        RECT  4.780 1.270 5.020 3.130 ;
        RECT  4.380 1.270 4.780 1.510 ;
        RECT  3.500 2.890 4.780 3.130 ;
        RECT  3.260 2.380 3.500 3.130 ;
        RECT  2.860 2.380 3.260 2.620 ;
        RECT  2.960 1.060 3.120 1.460 ;
        RECT  2.340 2.900 2.980 3.140 ;
        RECT  2.720 1.060 2.960 1.850 ;
        RECT  2.620 2.130 2.860 2.620 ;
        RECT  2.340 1.610 2.720 1.850 ;
        RECT  2.100 1.610 2.340 3.140 ;
        RECT  1.820 0.930 2.180 1.330 ;
        RECT  1.580 0.930 1.820 3.660 ;
        RECT  1.060 0.990 1.300 3.460 ;
    END
END MXI4X2

MACRO MXI4X1
    CLASS CORE ;
    FOREIGN MXI4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MXI4XL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.060 2.950 14.170 3.210 ;
        RECT  14.170 2.940 14.610 3.220 ;
        RECT  14.610 1.400 14.630 1.800 ;
        RECT  14.610 2.940 14.670 3.470 ;
        RECT  14.630 1.400 14.670 1.820 ;
        RECT  14.670 1.400 15.010 3.470 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  12.540 2.250 13.090 2.650 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.030 1.820 4.450 2.380 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.410 1.260 5.420 1.830 ;
        RECT  5.420 1.260 5.820 2.000 ;
        RECT  5.820 1.260 5.830 1.830 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.370 1.600 8.610 2.060 ;
        RECT  8.610 1.820 8.780 2.060 ;
        RECT  8.780 1.820 9.020 2.090 ;
        RECT  9.020 1.830 9.040 2.090 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.200 1.660 3.360 2.060 ;
        RECT  3.360 1.280 3.500 2.060 ;
        RECT  3.500 1.270 3.600 2.060 ;
        RECT  3.600 1.270 3.760 1.530 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.020 0.730 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 3.490 5.440 ;
        RECT  3.490 4.050 3.500 5.440 ;
        RECT  3.500 3.930 3.900 5.440 ;
        RECT  3.900 4.050 3.910 5.440 ;
        RECT  3.910 4.640 5.130 5.440 ;
        RECT  5.130 4.050 5.140 5.440 ;
        RECT  5.140 3.930 5.540 5.440 ;
        RECT  5.540 4.050 5.550 5.440 ;
        RECT  5.550 4.640 8.520 5.440 ;
        RECT  8.520 4.480 8.920 5.440 ;
        RECT  8.920 4.640 11.960 5.440 ;
        RECT  11.960 3.460 11.970 5.440 ;
        RECT  11.970 3.260 12.370 5.440 ;
        RECT  12.370 3.460 12.380 5.440 ;
        RECT  12.380 4.640 13.790 5.440 ;
        RECT  13.790 4.480 14.190 5.440 ;
        RECT  14.190 4.640 15.180 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.370 0.400 ;
        RECT  0.370 -0.400 0.770 0.560 ;
        RECT  0.770 -0.400 3.410 0.400 ;
        RECT  3.410 -0.400 3.420 0.870 ;
        RECT  3.420 -0.400 3.820 0.990 ;
        RECT  3.820 -0.400 3.830 0.870 ;
        RECT  3.830 -0.400 5.130 0.400 ;
        RECT  5.130 -0.400 5.140 0.870 ;
        RECT  5.140 -0.400 5.540 0.990 ;
        RECT  5.540 -0.400 5.550 0.870 ;
        RECT  5.550 -0.400 8.440 0.400 ;
        RECT  8.440 -0.400 8.840 0.560 ;
        RECT  8.840 -0.400 12.080 0.400 ;
        RECT  12.080 -0.400 12.090 0.750 ;
        RECT  12.090 -0.400 12.490 0.870 ;
        RECT  12.490 -0.400 12.500 0.750 ;
        RECT  12.500 -0.400 13.790 0.400 ;
        RECT  13.790 -0.400 14.190 0.560 ;
        RECT  14.190 -0.400 15.180 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.230 2.070 14.390 2.470 ;
        RECT  13.990 1.150 14.230 2.470 ;
        RECT  11.770 1.150 13.990 1.390 ;
        RECT  13.360 1.670 13.600 3.240 ;
        RECT  11.850 1.670 13.360 1.910 ;
        RECT  13.250 3.000 13.360 3.240 ;
        RECT  12.850 3.000 13.250 3.400 ;
        RECT  11.930 2.430 12.010 2.830 ;
        RECT  11.690 2.410 11.930 2.830 ;
        RECT  11.610 1.670 11.850 1.950 ;
        RECT  11.530 0.670 11.770 1.390 ;
        RECT  11.450 2.410 11.690 4.140 ;
        RECT  11.390 1.710 11.610 1.950 ;
        RECT  10.340 0.670 11.530 0.910 ;
        RECT  6.230 3.900 11.450 4.140 ;
        RECT  11.150 1.710 11.390 2.110 ;
        RECT  10.860 1.190 11.240 1.430 ;
        RECT  10.860 3.030 11.170 3.430 ;
        RECT  10.620 1.190 10.860 3.430 ;
        RECT  10.100 0.670 10.340 3.430 ;
        RECT  10.080 3.030 10.100 3.430 ;
        RECT  9.430 1.010 9.670 3.430 ;
        RECT  9.260 1.010 9.430 1.410 ;
        RECT  9.240 3.030 9.430 3.430 ;
        RECT  8.560 2.420 9.140 2.660 ;
        RECT  8.320 2.420 8.560 3.600 ;
        RECT  7.520 3.360 8.320 3.600 ;
        RECT  8.040 1.010 8.100 1.430 ;
        RECT  7.800 1.010 8.040 3.080 ;
        RECT  7.280 0.960 7.520 3.600 ;
        RECT  6.900 0.960 7.280 1.360 ;
        RECT  6.790 3.360 7.280 3.600 ;
        RECT  6.760 1.640 7.000 3.080 ;
        RECT  6.500 1.640 6.760 1.880 ;
        RECT  5.960 2.840 6.760 3.080 ;
        RECT  6.260 1.020 6.500 1.880 ;
        RECT  6.240 2.160 6.480 2.560 ;
        RECT  6.100 1.020 6.260 1.430 ;
        RECT  5.020 2.320 6.240 2.560 ;
        RECT  5.990 3.410 6.230 4.140 ;
        RECT  1.760 3.410 5.990 3.650 ;
        RECT  4.780 1.310 5.020 3.090 ;
        RECT  4.700 1.310 4.780 1.550 ;
        RECT  3.610 2.850 4.780 3.090 ;
        RECT  4.300 1.100 4.700 1.550 ;
        RECT  3.370 2.370 3.610 3.090 ;
        RECT  2.800 2.370 3.370 2.610 ;
        RECT  2.280 2.890 3.060 3.130 ;
        RECT  2.760 1.070 2.920 1.470 ;
        RECT  2.560 2.210 2.800 2.610 ;
        RECT  2.520 1.070 2.760 1.930 ;
        RECT  2.280 1.690 2.520 1.930 ;
        RECT  2.040 1.690 2.280 3.130 ;
        RECT  1.760 1.170 2.000 1.410 ;
        RECT  1.520 1.170 1.760 3.650 ;
        RECT  1.000 1.150 1.240 3.330 ;
        RECT  0.720 1.150 1.000 1.550 ;
    END
END MXI4X1

MACRO MXI2XL
    CLASS CORE ;
    FOREIGN MXI2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.710 1.190 2.950 3.410 ;
        RECT  2.950 2.390 3.090 3.410 ;
        RECT  3.090 2.390 3.100 2.650 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.740 2.170 1.140 2.660 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 1.830 1.490 2.110 ;
        RECT  1.490 1.830 1.890 2.360 ;
        RECT  1.890 1.830 1.900 2.110 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.970 2.010 4.160 2.470 ;
        RECT  4.160 1.830 4.420 2.470 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.040 5.440 ;
        RECT  1.040 4.060 1.050 5.440 ;
        RECT  1.050 3.940 1.450 5.440 ;
        RECT  1.450 4.060 1.460 5.440 ;
        RECT  1.460 4.640 4.060 5.440 ;
        RECT  4.060 4.480 4.460 5.440 ;
        RECT  4.460 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.080 0.400 ;
        RECT  1.080 -0.400 1.480 0.960 ;
        RECT  1.480 -0.400 4.060 0.400 ;
        RECT  4.060 -0.400 4.460 0.560 ;
        RECT  4.460 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.700 2.950 3.830 3.350 ;
        RECT  3.700 1.140 3.790 1.540 ;
        RECT  3.460 1.140 3.700 3.350 ;
        RECT  3.390 1.140 3.460 1.540 ;
        RECT  3.430 2.950 3.460 3.350 ;
        RECT  2.330 3.770 2.490 4.170 ;
        RECT  2.170 1.150 2.410 3.140 ;
        RECT  2.090 3.420 2.330 4.170 ;
        RECT  1.870 1.150 2.170 1.550 ;
        RECT  1.850 2.900 2.170 3.140 ;
        RECT  0.570 3.420 2.090 3.660 ;
        RECT  0.410 1.220 0.610 1.620 ;
        RECT  0.410 3.060 0.570 3.660 ;
        RECT  0.170 1.220 0.410 3.660 ;
    END
END MXI2XL

MACRO MXI2X4
    CLASS CORE ;
    FOREIGN MXI2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MXI2XL ;
    SIZE 9.900 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.500 0.680 4.070 1.080 ;
        RECT  2.820 3.540 4.360 3.780 ;
        RECT  4.070 0.680 4.360 2.410 ;
        RECT  4.360 0.680 4.510 3.780 ;
        RECT  4.510 1.980 4.640 3.780 ;
        RECT  4.510 0.680 4.870 0.980 ;
        RECT  4.640 3.500 4.950 3.780 ;
        RECT  4.870 0.680 5.690 0.920 ;
        RECT  5.690 0.680 6.170 1.080 ;
        RECT  4.950 3.540 6.270 3.780 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.300 3.940 2.540 4.360 ;
        RECT  2.540 4.060 2.970 4.360 ;
        RECT  2.970 4.120 5.610 4.360 ;
        RECT  5.610 4.050 6.530 4.370 ;
        RECT  6.530 2.870 6.550 4.370 ;
        RECT  6.550 2.870 6.770 4.360 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.030 2.160 8.510 2.660 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.710 2.180 0.860 2.580 ;
        RECT  0.860 2.180 1.120 2.650 ;
        RECT  1.120 2.180 1.690 2.580 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.230 0.170 5.440 ;
        RECT  0.170 4.030 0.570 5.440 ;
        RECT  0.570 4.230 0.580 5.440 ;
        RECT  0.580 4.640 1.730 5.440 ;
        RECT  1.730 4.020 1.970 5.440 ;
        RECT  1.970 4.640 7.620 5.440 ;
        RECT  7.620 3.870 7.630 5.440 ;
        RECT  7.630 3.670 8.030 5.440 ;
        RECT  8.030 3.870 8.040 5.440 ;
        RECT  8.040 4.640 9.140 5.440 ;
        RECT  9.140 4.220 9.150 5.440 ;
        RECT  9.150 4.020 9.550 5.440 ;
        RECT  9.550 4.220 9.560 5.440 ;
        RECT  9.560 4.640 9.900 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.360 0.400 ;
        RECT  0.360 -0.400 0.370 0.900 ;
        RECT  0.370 -0.400 0.770 1.100 ;
        RECT  0.770 -0.400 0.780 0.900 ;
        RECT  0.780 -0.400 1.640 0.400 ;
        RECT  1.640 -0.400 1.650 0.900 ;
        RECT  1.650 -0.400 2.050 1.100 ;
        RECT  2.050 -0.400 2.060 0.900 ;
        RECT  2.060 -0.400 7.680 0.400 ;
        RECT  7.680 -0.400 8.080 0.560 ;
        RECT  8.080 -0.400 9.010 0.400 ;
        RECT  9.010 -0.400 9.020 0.900 ;
        RECT  9.020 -0.400 9.420 1.100 ;
        RECT  9.420 -0.400 9.430 0.900 ;
        RECT  9.430 -0.400 9.900 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  9.030 1.540 9.270 3.170 ;
        RECT  8.750 1.540 9.030 1.780 ;
        RECT  8.820 2.930 9.030 3.170 ;
        RECT  8.420 2.930 8.820 3.330 ;
        RECT  8.590 1.380 8.750 1.780 ;
        RECT  8.350 0.860 8.590 1.780 ;
        RECT  6.690 0.860 8.350 1.100 ;
        RECT  7.210 2.250 7.350 3.150 ;
        RECT  7.110 1.380 7.210 3.150 ;
        RECT  6.970 1.380 7.110 2.490 ;
        RECT  5.750 2.250 6.970 2.490 ;
        RECT  6.450 0.860 6.690 1.600 ;
        RECT  5.470 1.360 6.450 1.600 ;
        RECT  5.450 1.360 5.470 3.210 ;
        RECT  5.230 1.230 5.450 3.210 ;
        RECT  5.050 1.230 5.230 1.600 ;
        RECT  5.070 2.810 5.230 3.210 ;
        RECT  3.560 2.810 3.960 3.210 ;
        RECT  2.250 2.930 3.560 3.170 ;
        RECT  3.110 1.360 3.510 1.780 ;
        RECT  2.250 1.540 3.110 1.780 ;
        RECT  2.010 1.540 2.250 3.170 ;
        RECT  1.380 1.540 2.010 1.780 ;
        RECT  1.310 2.930 2.010 3.170 ;
        RECT  0.980 1.380 1.380 1.780 ;
        RECT  0.910 2.930 1.310 3.330 ;
    END
END MXI2X4

MACRO MXI2X2
    CLASS CORE ;
    FOREIGN MXI2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MXI2XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.660 3.490 3.090 3.890 ;
        RECT  3.090 3.490 3.100 3.770 ;
        RECT  3.100 3.490 3.130 3.730 ;
        RECT  3.130 1.200 3.370 3.730 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.770 2.790 1.010 3.210 ;
        RECT  1.010 2.970 1.520 3.210 ;
        RECT  1.520 2.950 1.780 3.210 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 1.120 2.090 ;
        RECT  1.120 1.850 1.170 2.090 ;
        RECT  1.170 1.850 1.410 2.460 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.690 1.830 5.090 2.440 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.040 5.440 ;
        RECT  1.040 4.110 1.050 5.440 ;
        RECT  1.050 3.910 1.450 5.440 ;
        RECT  1.450 4.110 1.460 5.440 ;
        RECT  1.460 4.640 4.520 5.440 ;
        RECT  4.520 4.080 4.530 5.440 ;
        RECT  4.530 3.590 4.930 5.440 ;
        RECT  4.930 4.080 4.940 5.440 ;
        RECT  4.940 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        RECT  0.980 -0.400 0.990 0.830 ;
        RECT  0.990 -0.400 1.390 1.030 ;
        RECT  1.390 -0.400 1.400 0.830 ;
        RECT  1.400 -0.400 4.720 0.400 ;
        RECT  4.720 -0.400 5.120 0.560 ;
        RECT  5.120 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.170 1.380 4.410 3.310 ;
        RECT  4.050 3.070 4.170 3.310 ;
        RECT  3.650 3.070 4.050 4.050 ;
        RECT  3.650 0.680 3.890 2.430 ;
        RECT  1.930 0.680 3.650 0.920 ;
        RECT  2.610 1.500 2.850 3.210 ;
        RECT  2.210 1.340 2.610 1.740 ;
        RECT  2.380 2.970 2.610 3.210 ;
        RECT  2.140 2.970 2.380 4.230 ;
        RECT  1.930 2.250 2.330 2.650 ;
        RECT  1.810 3.830 2.140 4.230 ;
        RECT  1.690 0.680 1.930 2.650 ;
        RECT  0.570 1.310 1.690 1.550 ;
        RECT  0.450 3.480 0.630 3.880 ;
        RECT  0.450 1.050 0.570 1.550 ;
        RECT  0.230 1.050 0.450 3.880 ;
        RECT  0.210 1.050 0.230 3.860 ;
        RECT  0.170 1.050 0.210 1.450 ;
    END
END MXI2X2

MACRO MXI2X1
    CLASS CORE ;
    FOREIGN MXI2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MXI2XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.710 1.190 2.950 3.410 ;
        RECT  2.950 2.390 3.090 3.410 ;
        RECT  3.090 2.390 3.100 2.650 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.740 2.170 1.140 2.660 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 1.830 1.490 2.110 ;
        RECT  1.490 1.830 1.890 2.360 ;
        RECT  1.890 1.830 1.900 2.110 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.970 2.030 4.160 2.490 ;
        RECT  4.160 1.830 4.420 2.490 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.980 5.440 ;
        RECT  0.980 4.060 0.990 5.440 ;
        RECT  0.990 3.940 1.390 5.440 ;
        RECT  1.390 4.060 1.400 5.440 ;
        RECT  1.400 4.640 4.060 5.440 ;
        RECT  4.060 4.480 4.460 5.440 ;
        RECT  4.460 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.080 0.400 ;
        RECT  1.080 -0.400 1.090 1.270 ;
        RECT  1.090 -0.400 1.490 1.470 ;
        RECT  1.490 -0.400 1.500 1.270 ;
        RECT  1.500 -0.400 4.060 0.400 ;
        RECT  4.060 -0.400 4.460 0.560 ;
        RECT  4.460 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.700 2.950 3.830 3.350 ;
        RECT  3.700 1.140 3.790 1.540 ;
        RECT  3.460 1.140 3.700 3.350 ;
        RECT  3.390 1.140 3.460 1.540 ;
        RECT  3.430 2.950 3.460 3.350 ;
        RECT  2.330 3.920 2.490 4.320 ;
        RECT  2.170 1.150 2.410 3.140 ;
        RECT  2.090 3.420 2.330 4.320 ;
        RECT  1.870 1.150 2.170 1.550 ;
        RECT  1.850 2.900 2.170 3.140 ;
        RECT  0.570 3.420 2.090 3.660 ;
        RECT  0.410 1.220 0.610 1.620 ;
        RECT  0.410 3.060 0.570 3.660 ;
        RECT  0.170 1.220 0.410 3.660 ;
    END
END MXI2X1

MACRO MX4XL
    CLASS CORE ;
    FOREIGN MX4XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.630 2.940 12.690 4.340 ;
        RECT  12.690 1.390 12.930 4.340 ;
        RECT  12.930 1.470 12.990 4.340 ;
        RECT  12.990 2.940 13.030 4.340 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.100 0.660 9.700 0.980 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.110 2.210 4.530 2.660 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.280 1.660 3.500 2.080 ;
        RECT  3.500 1.660 3.680 2.090 ;
        RECT  3.680 1.830 3.760 2.090 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.460 2.500 ;
        RECT  0.460 1.900 0.800 2.500 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.400 1.270 5.820 2.020 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.280 1.870 8.290 2.270 ;
        RECT  8.290 1.840 8.780 2.270 ;
        RECT  8.780 1.830 9.040 2.270 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 3.610 5.440 ;
        RECT  3.610 4.110 3.620 5.440 ;
        RECT  3.620 3.990 4.020 5.440 ;
        RECT  4.020 4.110 4.030 5.440 ;
        RECT  4.030 4.640 5.230 5.440 ;
        RECT  5.230 4.110 5.240 5.440 ;
        RECT  5.240 3.990 5.640 5.440 ;
        RECT  5.640 4.110 5.650 5.440 ;
        RECT  5.650 4.640 8.500 5.440 ;
        RECT  8.500 4.480 8.900 5.440 ;
        RECT  8.900 4.640 11.810 5.440 ;
        RECT  11.810 4.480 12.210 5.440 ;
        RECT  12.210 4.640 13.200 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 3.450 0.400 ;
        RECT  3.450 -0.400 3.460 1.180 ;
        RECT  3.460 -0.400 3.860 1.380 ;
        RECT  3.860 -0.400 3.870 1.180 ;
        RECT  3.870 -0.400 5.270 0.400 ;
        RECT  5.270 -0.400 5.670 0.980 ;
        RECT  5.670 -0.400 8.370 0.400 ;
        RECT  8.370 -0.400 8.770 0.560 ;
        RECT  8.770 -0.400 12.440 0.400 ;
        RECT  12.440 -0.400 12.840 0.560 ;
        RECT  12.840 -0.400 13.200 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.170 0.860 12.410 2.360 ;
        RECT  11.150 0.860 12.170 1.100 ;
        RECT  11.890 2.820 11.980 3.220 ;
        RECT  11.810 1.380 11.890 3.220 ;
        RECT  11.650 1.380 11.810 4.180 ;
        RECT  11.570 2.820 11.650 4.180 ;
        RECT  6.590 3.940 11.570 4.180 ;
        RECT  11.070 3.030 11.220 3.430 ;
        RECT  11.070 0.860 11.150 1.510 ;
        RECT  10.910 0.860 11.070 3.430 ;
        RECT  10.830 1.110 10.910 3.430 ;
        RECT  10.750 1.110 10.830 1.510 ;
        RECT  10.820 3.030 10.830 3.430 ;
        RECT  10.300 1.190 10.450 3.400 ;
        RECT  10.290 1.110 10.300 3.400 ;
        RECT  10.210 1.110 10.290 3.660 ;
        RECT  10.060 1.110 10.210 1.510 ;
        RECT  10.050 3.000 10.210 3.660 ;
        RECT  7.490 3.420 10.050 3.660 ;
        RECT  9.770 1.820 9.930 2.220 ;
        RECT  9.700 1.280 9.770 2.220 ;
        RECT  9.700 2.900 9.710 3.140 ;
        RECT  9.460 1.280 9.700 3.140 ;
        RECT  9.240 1.280 9.460 1.520 ;
        RECT  9.310 2.900 9.460 3.140 ;
        RECT  7.770 1.000 8.010 3.140 ;
        RECT  7.250 1.080 7.490 3.660 ;
        RECT  6.930 1.080 7.250 1.320 ;
        RECT  6.950 3.330 7.250 3.660 ;
        RECT  6.730 1.610 6.970 3.050 ;
        RECT  6.870 3.330 6.950 3.570 ;
        RECT  6.570 1.610 6.730 1.850 ;
        RECT  6.510 2.810 6.730 3.050 ;
        RECT  6.350 3.470 6.590 4.180 ;
        RECT  6.330 1.000 6.570 1.850 ;
        RECT  6.110 2.810 6.510 3.190 ;
        RECT  6.210 2.130 6.450 2.530 ;
        RECT  2.200 3.470 6.350 3.710 ;
        RECT  6.170 1.000 6.330 1.400 ;
        RECT  5.040 2.290 6.210 2.530 ;
        RECT  4.800 1.410 5.040 3.170 ;
        RECT  4.740 1.410 4.800 1.650 ;
        RECT  3.590 2.930 4.800 3.170 ;
        RECT  4.340 1.250 4.740 1.650 ;
        RECT  3.350 2.370 3.590 3.170 ;
        RECT  2.880 2.370 3.350 2.610 ;
        RECT  2.360 2.890 3.040 3.130 ;
        RECT  2.820 1.060 2.980 1.460 ;
        RECT  2.640 2.210 2.880 2.610 ;
        RECT  2.580 1.060 2.820 1.850 ;
        RECT  2.360 1.610 2.580 1.850 ;
        RECT  2.120 1.610 2.360 3.130 ;
        RECT  1.840 1.090 2.200 1.330 ;
        RECT  1.880 3.410 2.200 3.710 ;
        RECT  1.840 3.410 1.880 3.650 ;
        RECT  1.600 1.090 1.840 3.650 ;
        RECT  1.080 1.040 1.320 3.460 ;
    END
END MX4XL

MACRO MX4X4
    CLASS CORE ;
    FOREIGN MX4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MX4XL ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.630 1.820 14.650 3.220 ;
        RECT  14.650 1.350 14.660 3.220 ;
        RECT  14.660 1.150 15.060 3.720 ;
        RECT  15.060 1.350 15.070 3.220 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  10.890 2.300 11.130 3.780 ;
        RECT  11.130 2.300 11.290 2.540 ;
        RECT  11.130 3.500 12.950 3.780 ;
        RECT  12.950 2.380 13.190 3.780 ;
        RECT  13.190 3.500 13.200 3.780 ;
        RECT  13.190 2.380 13.510 2.790 ;
        RECT  13.510 2.390 13.590 2.790 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.020 4.080 2.180 4.320 ;
        RECT  2.180 4.070 2.440 4.330 ;
        RECT  2.440 4.080 2.850 4.320 ;
        RECT  2.850 3.940 3.090 4.320 ;
        RECT  3.090 3.940 5.190 4.180 ;
        RECT  5.190 3.890 5.590 4.180 ;
        RECT  5.590 3.940 7.640 4.180 ;
        RECT  7.640 3.940 7.880 4.370 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.720 2.190 3.960 2.590 ;
        RECT  3.960 2.350 4.160 2.590 ;
        RECT  4.160 2.350 4.410 2.650 ;
        RECT  4.410 2.390 4.420 2.650 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.210 2.090 ;
        RECT  0.210 1.830 0.460 2.460 ;
        RECT  0.460 1.840 0.730 2.460 ;
        RECT  0.730 1.840 0.810 2.240 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.960 1.750 6.490 2.110 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.220 2.200 9.360 2.600 ;
        RECT  9.360 2.200 9.440 2.640 ;
        RECT  9.440 2.200 9.620 2.650 ;
        RECT  9.620 2.390 9.700 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.000 0.170 5.440 ;
        RECT  0.170 3.510 0.570 5.440 ;
        RECT  0.570 4.000 0.580 5.440 ;
        RECT  0.580 4.640 3.930 5.440 ;
        RECT  3.930 4.480 4.330 5.440 ;
        RECT  4.330 4.640 5.650 5.440 ;
        RECT  5.650 4.480 6.050 5.440 ;
        RECT  6.050 4.640 9.500 5.440 ;
        RECT  9.500 4.480 9.900 5.440 ;
        RECT  9.900 4.640 13.980 5.440 ;
        RECT  13.980 4.230 13.990 5.440 ;
        RECT  13.990 4.030 14.390 5.440 ;
        RECT  14.390 4.230 14.400 5.440 ;
        RECT  14.400 4.640 15.260 5.440 ;
        RECT  15.260 4.230 15.270 5.440 ;
        RECT  15.270 4.030 15.670 5.440 ;
        RECT  15.670 4.230 15.680 5.440 ;
        RECT  15.680 4.640 15.840 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 0.790 ;
        RECT  0.170 -0.400 0.570 0.990 ;
        RECT  0.570 -0.400 0.580 0.790 ;
        RECT  0.580 -0.400 3.930 0.400 ;
        RECT  3.930 -0.400 4.330 0.560 ;
        RECT  4.330 -0.400 5.680 0.400 ;
        RECT  5.680 -0.400 6.080 0.560 ;
        RECT  6.080 -0.400 9.500 0.400 ;
        RECT  9.500 -0.400 9.900 0.560 ;
        RECT  9.900 -0.400 13.980 0.400 ;
        RECT  13.980 -0.400 13.990 0.670 ;
        RECT  13.990 -0.400 14.390 0.870 ;
        RECT  14.390 -0.400 14.400 0.670 ;
        RECT  14.400 -0.400 15.260 0.400 ;
        RECT  15.260 -0.400 15.270 0.670 ;
        RECT  15.270 -0.400 15.670 0.870 ;
        RECT  15.670 -0.400 15.680 0.670 ;
        RECT  15.680 -0.400 15.840 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.090 1.150 14.330 3.310 ;
        RECT  13.430 1.150 14.090 1.390 ;
        RECT  13.710 3.070 14.090 3.310 ;
        RECT  12.680 1.670 13.810 2.070 ;
        RECT  13.470 3.070 13.710 4.290 ;
        RECT  10.610 4.050 13.470 4.290 ;
        RECT  13.030 0.970 13.430 1.390 ;
        RECT  12.670 1.330 12.680 2.070 ;
        RECT  12.490 0.980 12.670 2.070 ;
        RECT  12.250 0.980 12.490 3.230 ;
        RECT  12.090 2.830 12.250 3.230 ;
        RECT  11.810 0.810 11.910 1.210 ;
        RECT  11.570 0.810 11.810 3.230 ;
        RECT  11.510 0.810 11.570 1.210 ;
        RECT  11.410 2.830 11.570 3.230 ;
        RECT  8.320 0.860 11.510 1.100 ;
        RECT  10.690 1.490 11.290 1.890 ;
        RECT  10.610 1.380 10.690 1.890 ;
        RECT  10.370 1.380 10.610 3.360 ;
        RECT  10.370 3.940 10.610 4.290 ;
        RECT  10.290 1.380 10.370 1.620 ;
        RECT  8.400 3.940 10.370 4.180 ;
        RECT  8.920 1.380 9.080 1.620 ;
        RECT  8.920 3.260 9.080 3.660 ;
        RECT  8.680 1.380 8.920 3.660 ;
        RECT  8.160 3.420 8.400 4.180 ;
        RECT  8.130 0.860 8.320 1.330 ;
        RECT  8.130 2.900 8.290 3.140 ;
        RECT  6.190 3.420 8.160 3.660 ;
        RECT  7.890 0.860 8.130 3.140 ;
        RECT  7.370 1.190 7.610 3.140 ;
        RECT  7.160 1.190 7.370 1.590 ;
        RECT  6.470 2.900 7.370 3.140 ;
        RECT  6.880 0.670 7.230 0.910 ;
        RECT  6.850 1.940 7.090 2.620 ;
        RECT  6.640 0.670 6.880 1.100 ;
        RECT  5.180 2.380 6.850 2.620 ;
        RECT  3.380 0.860 6.640 1.100 ;
        RECT  5.950 3.370 6.190 3.660 ;
        RECT  4.820 3.370 5.950 3.610 ;
        RECT  5.090 2.380 5.180 3.090 ;
        RECT  4.780 1.450 5.090 3.090 ;
        RECT  4.580 3.370 4.820 3.660 ;
        RECT  3.370 1.450 4.780 1.690 ;
        RECT  2.090 3.420 4.580 3.660 ;
        RECT  2.460 2.900 3.510 3.140 ;
        RECT  3.140 0.670 3.380 1.100 ;
        RECT  3.130 1.450 3.370 2.570 ;
        RECT  2.780 0.670 3.140 0.910 ;
        RECT  2.740 2.170 3.130 2.570 ;
        RECT  2.460 1.230 2.850 1.630 ;
        RECT  2.450 1.230 2.460 3.140 ;
        RECT  2.220 1.390 2.450 3.140 ;
        RECT  1.930 0.710 2.090 1.110 ;
        RECT  1.930 3.420 2.090 3.710 ;
        RECT  1.690 0.710 1.930 3.710 ;
        RECT  1.090 0.930 1.330 4.200 ;
        RECT  0.930 0.930 1.090 1.330 ;
        RECT  0.930 3.220 1.090 4.200 ;
    END
END MX4X4

MACRO MX4X2
    CLASS CORE ;
    FOREIGN MX4X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MX4XL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.600 3.700 14.610 4.160 ;
        RECT  14.610 2.940 14.690 4.160 ;
        RECT  14.610 0.960 14.690 1.360 ;
        RECT  14.690 0.960 14.930 4.160 ;
        RECT  14.930 2.940 15.010 4.160 ;
        RECT  14.930 0.960 15.010 1.360 ;
        RECT  15.010 3.700 15.020 4.160 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  10.880 3.500 10.890 3.780 ;
        RECT  10.890 2.300 11.130 3.780 ;
        RECT  11.130 2.300 11.290 2.540 ;
        RECT  11.130 3.500 12.810 3.780 ;
        RECT  12.810 2.380 13.050 3.780 ;
        RECT  13.050 3.500 13.060 3.780 ;
        RECT  13.050 2.380 13.510 2.790 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.020 4.080 2.180 4.320 ;
        RECT  2.180 4.070 2.440 4.330 ;
        RECT  2.440 4.080 2.850 4.320 ;
        RECT  2.850 3.940 3.090 4.320 ;
        RECT  3.090 3.940 5.190 4.180 ;
        RECT  5.190 3.890 5.590 4.180 ;
        RECT  5.590 3.940 7.640 4.180 ;
        RECT  7.640 3.940 7.880 4.370 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.720 2.190 3.960 2.590 ;
        RECT  3.960 2.350 4.160 2.590 ;
        RECT  4.160 2.350 4.410 2.650 ;
        RECT  4.410 2.390 4.420 2.650 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.460 2.480 ;
        RECT  0.460 1.840 0.550 2.480 ;
        RECT  0.550 1.840 0.810 2.240 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.960 1.750 6.490 2.110 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.220 2.200 9.360 2.600 ;
        RECT  9.360 2.200 9.440 2.640 ;
        RECT  9.440 2.200 9.620 2.650 ;
        RECT  9.620 2.390 9.700 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.000 0.170 5.440 ;
        RECT  0.170 3.510 0.570 5.440 ;
        RECT  0.570 4.000 0.580 5.440 ;
        RECT  0.580 4.640 3.930 5.440 ;
        RECT  3.930 4.480 4.330 5.440 ;
        RECT  4.330 4.640 5.650 5.440 ;
        RECT  5.650 4.480 6.050 5.440 ;
        RECT  6.050 4.640 9.500 5.440 ;
        RECT  9.500 4.480 9.900 5.440 ;
        RECT  9.900 4.640 13.840 5.440 ;
        RECT  13.840 4.130 13.850 5.440 ;
        RECT  13.850 3.930 14.250 5.440 ;
        RECT  14.250 4.130 14.260 5.440 ;
        RECT  14.260 4.640 15.180 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 0.790 ;
        RECT  0.170 -0.400 0.570 0.990 ;
        RECT  0.570 -0.400 0.580 0.790 ;
        RECT  0.580 -0.400 3.930 0.400 ;
        RECT  3.930 -0.400 4.330 0.560 ;
        RECT  4.330 -0.400 5.680 0.400 ;
        RECT  5.680 -0.400 6.080 0.560 ;
        RECT  6.080 -0.400 9.500 0.400 ;
        RECT  9.500 -0.400 9.900 0.560 ;
        RECT  9.900 -0.400 13.840 0.400 ;
        RECT  13.840 -0.400 13.850 0.670 ;
        RECT  13.850 -0.400 14.250 0.870 ;
        RECT  14.250 -0.400 14.260 0.670 ;
        RECT  14.260 -0.400 15.180 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.090 1.150 14.330 3.310 ;
        RECT  13.430 1.150 14.090 1.390 ;
        RECT  13.570 3.070 14.090 3.310 ;
        RECT  12.680 1.670 13.810 2.070 ;
        RECT  13.330 3.070 13.570 4.290 ;
        RECT  13.030 0.970 13.430 1.390 ;
        RECT  10.610 4.050 13.330 4.290 ;
        RECT  12.670 1.330 12.680 2.070 ;
        RECT  12.490 0.980 12.670 2.070 ;
        RECT  12.250 0.980 12.490 3.230 ;
        RECT  12.090 2.830 12.250 3.230 ;
        RECT  11.810 0.810 11.910 1.210 ;
        RECT  11.570 0.810 11.810 3.230 ;
        RECT  11.510 0.810 11.570 1.210 ;
        RECT  11.410 2.830 11.570 3.230 ;
        RECT  8.320 0.860 11.510 1.100 ;
        RECT  10.690 1.490 11.290 1.890 ;
        RECT  10.610 1.380 10.690 1.890 ;
        RECT  10.370 1.380 10.610 3.360 ;
        RECT  10.370 3.940 10.610 4.290 ;
        RECT  10.290 1.380 10.370 1.620 ;
        RECT  8.400 3.940 10.370 4.180 ;
        RECT  8.920 1.380 9.080 1.620 ;
        RECT  8.920 3.260 9.080 3.660 ;
        RECT  8.680 1.380 8.920 3.660 ;
        RECT  8.160 3.420 8.400 4.180 ;
        RECT  8.130 0.860 8.320 1.330 ;
        RECT  8.130 2.900 8.290 3.140 ;
        RECT  6.190 3.420 8.160 3.660 ;
        RECT  7.890 0.860 8.130 3.140 ;
        RECT  7.370 1.190 7.610 3.140 ;
        RECT  7.160 1.190 7.370 1.590 ;
        RECT  6.470 2.900 7.370 3.140 ;
        RECT  6.880 0.670 7.230 0.910 ;
        RECT  6.850 1.940 7.090 2.620 ;
        RECT  6.640 0.670 6.880 1.100 ;
        RECT  5.180 2.380 6.850 2.620 ;
        RECT  3.380 0.860 6.640 1.100 ;
        RECT  5.950 3.370 6.190 3.660 ;
        RECT  4.820 3.370 5.950 3.610 ;
        RECT  5.090 2.380 5.180 3.090 ;
        RECT  4.780 1.450 5.090 3.090 ;
        RECT  4.580 3.370 4.820 3.660 ;
        RECT  3.370 1.450 4.780 1.690 ;
        RECT  2.090 3.420 4.580 3.660 ;
        RECT  2.460 2.900 3.510 3.140 ;
        RECT  3.140 0.670 3.380 1.100 ;
        RECT  3.130 1.450 3.370 2.570 ;
        RECT  2.780 0.670 3.140 0.910 ;
        RECT  2.740 2.170 3.130 2.570 ;
        RECT  2.460 1.230 2.850 1.630 ;
        RECT  2.450 1.230 2.460 3.140 ;
        RECT  2.220 1.390 2.450 3.140 ;
        RECT  1.930 0.710 2.090 1.110 ;
        RECT  1.930 3.420 2.090 3.710 ;
        RECT  1.690 0.710 1.930 3.710 ;
        RECT  1.090 0.930 1.330 4.200 ;
        RECT  0.930 0.930 1.090 1.330 ;
        RECT  0.930 3.220 1.090 4.200 ;
    END
END MX4X2

MACRO MX4X1
    CLASS CORE ;
    FOREIGN MX4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MX4XL ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.630 3.750 12.710 4.150 ;
        RECT  12.710 0.670 12.990 4.150 ;
        RECT  12.990 2.950 13.000 3.210 ;
        RECT  12.990 3.750 13.030 4.150 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.180 0.660 9.780 0.980 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.110 2.210 4.530 2.660 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.280 1.740 3.680 2.140 ;
        RECT  3.680 1.830 3.760 2.090 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.210 2.090 ;
        RECT  0.210 1.830 0.460 2.460 ;
        RECT  0.460 2.060 0.800 2.460 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.400 1.270 5.410 2.020 ;
        RECT  5.410 1.270 5.810 2.060 ;
        RECT  5.810 1.270 5.820 2.020 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.280 1.870 8.290 2.270 ;
        RECT  8.290 1.840 8.780 2.270 ;
        RECT  8.780 1.830 9.040 2.270 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 3.610 5.440 ;
        RECT  3.610 4.110 3.620 5.440 ;
        RECT  3.620 3.990 4.020 5.440 ;
        RECT  4.020 4.110 4.030 5.440 ;
        RECT  4.030 4.640 5.100 5.440 ;
        RECT  5.100 4.110 5.110 5.440 ;
        RECT  5.110 3.990 5.510 5.440 ;
        RECT  5.510 4.110 5.520 5.440 ;
        RECT  5.520 4.640 8.500 5.440 ;
        RECT  8.500 4.480 8.900 5.440 ;
        RECT  8.900 4.640 11.810 5.440 ;
        RECT  11.810 4.480 12.210 5.440 ;
        RECT  12.210 4.640 13.200 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 3.390 0.400 ;
        RECT  3.390 -0.400 3.400 1.110 ;
        RECT  3.400 -0.400 3.800 1.310 ;
        RECT  3.800 -0.400 3.810 1.110 ;
        RECT  3.810 -0.400 5.260 0.400 ;
        RECT  5.260 -0.400 5.270 0.860 ;
        RECT  5.270 -0.400 5.670 0.980 ;
        RECT  5.670 -0.400 5.680 0.860 ;
        RECT  5.680 -0.400 8.510 0.400 ;
        RECT  8.510 -0.400 8.910 0.560 ;
        RECT  8.910 -0.400 11.810 0.400 ;
        RECT  11.810 -0.400 12.210 0.560 ;
        RECT  12.210 -0.400 13.200 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.170 0.860 12.410 2.390 ;
        RECT  11.150 0.860 12.170 1.100 ;
        RECT  11.890 2.820 11.980 3.220 ;
        RECT  11.810 1.410 11.890 3.220 ;
        RECT  11.650 1.410 11.810 4.180 ;
        RECT  11.570 2.820 11.650 4.180 ;
        RECT  6.590 3.940 11.570 4.180 ;
        RECT  11.150 3.030 11.220 3.430 ;
        RECT  10.910 0.860 11.150 3.430 ;
        RECT  10.750 1.110 10.910 1.510 ;
        RECT  10.820 3.030 10.910 3.430 ;
        RECT  10.370 3.260 10.450 3.660 ;
        RECT  10.130 1.100 10.370 3.660 ;
        RECT  10.060 1.100 10.130 1.500 ;
        RECT  10.050 3.260 10.130 3.660 ;
        RECT  7.490 3.420 10.050 3.660 ;
        RECT  9.780 1.780 9.810 2.180 ;
        RECT  9.720 1.280 9.780 2.180 ;
        RECT  9.710 1.280 9.720 2.930 ;
        RECT  9.410 1.280 9.710 3.140 ;
        RECT  9.240 1.280 9.410 1.520 ;
        RECT  9.310 2.900 9.410 3.140 ;
        RECT  7.770 1.050 8.010 3.140 ;
        RECT  7.250 1.080 7.490 3.660 ;
        RECT  6.930 1.080 7.250 1.320 ;
        RECT  6.870 3.420 7.250 3.660 ;
        RECT  6.730 1.610 6.970 3.140 ;
        RECT  6.520 1.610 6.730 1.850 ;
        RECT  6.510 2.900 6.730 3.140 ;
        RECT  6.350 3.470 6.590 4.180 ;
        RECT  6.280 1.000 6.520 1.850 ;
        RECT  6.110 2.900 6.510 3.190 ;
        RECT  6.210 2.170 6.450 2.580 ;
        RECT  2.200 3.470 6.350 3.710 ;
        RECT  6.120 1.000 6.280 1.400 ;
        RECT  5.040 2.340 6.210 2.580 ;
        RECT  4.800 1.410 5.040 3.190 ;
        RECT  4.680 1.410 4.800 1.650 ;
        RECT  3.590 2.950 4.800 3.190 ;
        RECT  4.280 1.110 4.680 1.650 ;
        RECT  3.350 2.420 3.590 3.190 ;
        RECT  2.880 2.420 3.350 2.660 ;
        RECT  2.360 2.950 3.040 3.190 ;
        RECT  2.820 1.060 2.980 1.460 ;
        RECT  2.640 2.210 2.880 2.660 ;
        RECT  2.580 1.060 2.820 1.850 ;
        RECT  2.360 1.610 2.580 1.850 ;
        RECT  2.120 1.610 2.360 3.190 ;
        RECT  1.840 1.090 2.200 1.330 ;
        RECT  1.840 3.470 2.200 3.870 ;
        RECT  1.600 1.090 1.840 3.870 ;
        RECT  1.080 1.040 1.320 3.460 ;
    END
END MX4X1

MACRO MX2XL
    CLASS CORE ;
    FOREIGN MX2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.820 1.270 4.930 1.530 ;
        RECT  4.930 1.260 5.250 1.540 ;
        RECT  5.190 3.310 5.350 3.710 ;
        RECT  5.250 1.080 5.350 1.540 ;
        RECT  5.350 1.080 5.590 3.710 ;
        RECT  5.590 1.080 5.650 1.480 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.740 1.820 1.210 2.240 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.190 2.660 1.230 3.200 ;
        RECT  1.230 2.650 1.520 3.200 ;
        RECT  1.520 2.650 1.600 3.210 ;
        RECT  1.600 2.950 1.780 3.210 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.050 1.820 4.510 2.260 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.040 5.440 ;
        RECT  1.040 3.690 1.050 5.440 ;
        RECT  1.050 3.490 1.450 5.440 ;
        RECT  1.450 3.690 1.460 5.440 ;
        RECT  1.460 4.640 4.360 5.440 ;
        RECT  4.360 4.480 4.760 5.440 ;
        RECT  4.760 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.040 0.400 ;
        RECT  1.040 -0.400 1.050 0.830 ;
        RECT  1.050 -0.400 1.450 1.030 ;
        RECT  1.450 -0.400 1.460 0.830 ;
        RECT  1.460 -0.400 4.360 0.400 ;
        RECT  4.360 -0.400 4.760 0.560 ;
        RECT  4.760 -0.400 5.940 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.890 2.550 5.050 2.950 ;
        RECT  4.650 2.550 4.890 4.070 ;
        RECT  3.280 3.830 4.650 4.070 ;
        RECT  3.560 1.000 3.800 3.550 ;
        RECT  3.040 1.070 3.280 4.070 ;
        RECT  2.690 1.070 3.040 1.310 ;
        RECT  2.690 3.310 3.040 3.710 ;
        RECT  2.520 1.590 2.760 3.030 ;
        RECT  2.250 1.590 2.520 1.830 ;
        RECT  2.390 2.790 2.520 3.030 ;
        RECT  2.150 2.790 2.390 3.730 ;
        RECT  2.010 1.000 2.250 1.830 ;
        RECT  1.990 2.110 2.230 2.510 ;
        RECT  1.930 3.490 2.150 3.730 ;
        RECT  1.720 2.110 1.990 2.350 ;
        RECT  1.480 1.310 1.720 2.350 ;
        RECT  0.570 1.310 1.480 1.550 ;
        RECT  0.410 1.130 0.570 1.550 ;
        RECT  0.410 3.110 0.570 3.510 ;
        RECT  0.170 1.130 0.410 3.510 ;
    END
END MX2XL

MACRO MX2X4
    CLASS CORE ;
    FOREIGN MX2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MX2XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  5.210 3.940 5.610 4.370 ;
        RECT  5.390 0.700 5.830 2.100 ;
        RECT  5.610 3.940 6.050 4.180 ;
        RECT  6.050 3.620 6.060 4.180 ;
        RECT  5.830 1.820 6.060 2.100 ;
        RECT  6.060 1.820 6.300 4.180 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.890 0.920 3.290 ;
        RECT  0.920 2.960 1.520 3.200 ;
        RECT  1.520 2.950 1.780 3.210 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.680 1.450 2.090 ;
        RECT  1.450 1.680 1.460 2.050 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 1.800 4.580 2.220 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.920 5.440 ;
        RECT  0.920 3.770 0.930 5.440 ;
        RECT  0.930 3.570 1.330 5.440 ;
        RECT  1.330 3.770 1.340 5.440 ;
        RECT  1.340 4.640 4.440 5.440 ;
        RECT  4.440 4.330 4.450 5.440 ;
        RECT  4.450 4.130 4.850 5.440 ;
        RECT  4.850 4.330 4.860 5.440 ;
        RECT  4.860 4.640 6.030 5.440 ;
        RECT  6.030 4.480 6.430 5.440 ;
        RECT  6.430 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.920 0.400 ;
        RECT  0.920 -0.400 0.930 1.190 ;
        RECT  0.930 -0.400 1.330 1.390 ;
        RECT  1.330 -0.400 1.340 1.190 ;
        RECT  1.340 -0.400 4.650 0.400 ;
        RECT  4.650 -0.400 5.070 0.920 ;
        RECT  5.070 -0.400 6.100 0.400 ;
        RECT  6.100 -0.400 6.340 0.910 ;
        RECT  6.340 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.620 2.370 5.780 2.610 ;
        RECT  5.380 2.370 5.620 3.270 ;
        RECT  4.450 3.030 5.380 3.270 ;
        RECT  4.850 1.270 5.090 2.740 ;
        RECT  4.070 1.270 4.850 1.510 ;
        RECT  3.930 2.500 4.850 2.740 ;
        RECT  4.210 3.030 4.450 3.830 ;
        RECT  3.250 3.590 4.210 3.830 ;
        RECT  3.690 2.500 3.930 3.310 ;
        RECT  3.530 0.670 3.770 2.180 ;
        RECT  3.530 2.910 3.690 3.310 ;
        RECT  1.970 0.670 3.530 0.910 ;
        RECT  3.010 1.190 3.250 3.870 ;
        RECT  2.660 3.470 3.010 3.870 ;
        RECT  2.490 1.190 2.730 3.190 ;
        RECT  2.250 1.190 2.490 1.590 ;
        RECT  2.380 2.950 2.490 3.190 ;
        RECT  2.140 2.950 2.380 3.750 ;
        RECT  1.970 1.920 2.210 2.320 ;
        RECT  2.090 3.510 2.140 3.750 ;
        RECT  1.690 3.510 2.090 3.910 ;
        RECT  1.730 0.670 1.970 2.610 ;
        RECT  0.430 2.370 1.730 2.610 ;
        RECT  0.430 1.000 0.570 1.400 ;
        RECT  0.400 3.590 0.570 3.990 ;
        RECT  0.400 1.000 0.430 2.610 ;
        RECT  0.160 1.000 0.400 3.990 ;
    END
END MX2X4

MACRO MX2X2
    CLASS CORE ;
    FOREIGN MX2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MX2XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  5.360 3.210 5.480 4.190 ;
        RECT  5.480 2.950 5.540 4.190 ;
        RECT  5.440 0.870 5.540 1.400 ;
        RECT  5.540 0.870 5.760 4.190 ;
        RECT  5.760 0.870 5.780 4.180 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.750 2.810 1.150 3.210 ;
        RECT  1.150 2.960 1.520 3.200 ;
        RECT  1.520 2.950 1.780 3.210 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 1.120 2.090 ;
        RECT  1.120 1.850 1.200 2.090 ;
        RECT  1.200 1.850 1.440 2.370 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.300 1.300 4.540 2.120 ;
        RECT  4.540 1.300 4.820 1.540 ;
        RECT  4.820 1.270 5.060 1.540 ;
        RECT  5.060 1.270 5.080 1.530 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.130 5.440 ;
        RECT  1.130 3.690 1.140 5.440 ;
        RECT  1.140 3.490 1.540 5.440 ;
        RECT  1.540 3.690 1.550 5.440 ;
        RECT  1.550 4.640 4.540 5.440 ;
        RECT  4.540 4.480 4.940 5.440 ;
        RECT  4.940 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.150 0.400 ;
        RECT  1.150 -0.400 1.160 0.830 ;
        RECT  1.160 -0.400 1.560 1.030 ;
        RECT  1.560 -0.400 1.570 0.830 ;
        RECT  1.570 -0.400 4.580 0.400 ;
        RECT  4.580 -0.400 4.590 0.790 ;
        RECT  4.590 -0.400 4.990 0.990 ;
        RECT  4.990 -0.400 5.000 0.790 ;
        RECT  5.000 -0.400 5.940 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.020 1.960 5.260 2.670 ;
        RECT  4.540 2.430 5.020 2.670 ;
        RECT  4.300 2.430 4.540 4.180 ;
        RECT  3.500 3.940 4.300 4.180 ;
        RECT  3.780 1.000 4.020 3.670 ;
        RECT  3.260 1.140 3.500 4.180 ;
        RECT  3.180 1.140 3.260 1.380 ;
        RECT  2.830 3.480 3.260 3.880 ;
        RECT  2.780 0.980 3.180 1.380 ;
        RECT  2.740 1.660 2.980 3.200 ;
        RECT  2.480 1.660 2.740 1.900 ;
        RECT  2.400 2.960 2.740 3.200 ;
        RECT  2.240 0.790 2.480 1.900 ;
        RECT  2.230 2.180 2.470 2.620 ;
        RECT  2.390 2.960 2.400 3.560 ;
        RECT  2.150 2.950 2.390 3.930 ;
        RECT  2.040 0.790 2.240 1.030 ;
        RECT  1.960 2.180 2.230 2.420 ;
        RECT  1.720 1.310 1.960 2.420 ;
        RECT  0.570 1.310 1.720 1.550 ;
        RECT  0.470 3.490 0.630 3.890 ;
        RECT  0.470 1.040 0.570 1.550 ;
        RECT  0.230 1.040 0.470 3.890 ;
        RECT  0.170 1.040 0.230 1.440 ;
    END
END MX2X2

MACRO MX2X1
    CLASS CORE ;
    FOREIGN MX2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ MX2XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.820 1.270 4.930 1.530 ;
        RECT  4.930 1.260 5.180 1.540 ;
        RECT  5.180 3.310 5.340 3.710 ;
        RECT  5.180 1.120 5.340 1.540 ;
        RECT  5.340 1.120 5.580 3.710 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.750 1.820 1.210 2.240 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.190 2.660 1.230 3.200 ;
        RECT  1.230 2.650 1.520 3.200 ;
        RECT  1.520 2.650 1.600 3.210 ;
        RECT  1.600 2.950 1.780 3.210 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.030 1.820 4.510 2.240 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.090 5.440 ;
        RECT  1.090 3.610 1.100 5.440 ;
        RECT  1.100 3.490 1.500 5.440 ;
        RECT  1.500 3.610 1.510 5.440 ;
        RECT  1.510 4.640 4.320 5.440 ;
        RECT  4.320 4.480 4.720 5.440 ;
        RECT  4.720 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.040 0.400 ;
        RECT  1.040 -0.400 1.050 0.830 ;
        RECT  1.050 -0.400 1.450 1.030 ;
        RECT  1.450 -0.400 1.460 0.830 ;
        RECT  1.460 -0.400 4.290 0.400 ;
        RECT  4.290 -0.400 4.690 0.560 ;
        RECT  4.690 -0.400 5.940 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.890 2.580 5.060 2.980 ;
        RECT  4.650 2.580 4.890 4.070 ;
        RECT  3.270 3.830 4.650 4.070 ;
        RECT  3.550 1.000 3.790 3.550 ;
        RECT  3.030 1.070 3.270 4.070 ;
        RECT  2.690 1.070 3.030 1.310 ;
        RECT  2.700 3.310 3.030 3.710 ;
        RECT  2.510 1.590 2.750 3.030 ;
        RECT  2.240 1.590 2.510 1.830 ;
        RECT  2.380 2.790 2.510 3.030 ;
        RECT  2.140 2.790 2.380 3.730 ;
        RECT  2.000 1.000 2.240 1.830 ;
        RECT  1.990 2.110 2.230 2.510 ;
        RECT  1.860 3.490 2.140 3.730 ;
        RECT  1.720 2.110 1.990 2.350 ;
        RECT  1.480 1.310 1.720 2.350 ;
        RECT  0.570 1.310 1.480 1.550 ;
        RECT  0.410 1.090 0.570 1.550 ;
        RECT  0.410 3.110 0.570 3.510 ;
        RECT  0.170 1.090 0.410 3.510 ;
    END
END MX2X1

MACRO JKFFSRXL
    CLASS CORE ;
    FOREIGN JKFFSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.440 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.370 2.230 7.830 2.660 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.440 1.270 9.550 1.530 ;
        RECT  9.550 1.270 9.700 1.950 ;
        RECT  9.700 1.280 9.790 1.950 ;
        RECT  9.790 1.710 10.160 1.950 ;
        RECT  10.160 1.710 10.400 2.120 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  20.130 0.670 20.530 1.100 ;
        RECT  20.490 3.520 20.660 4.220 ;
        RECT  20.660 3.510 20.730 4.220 ;
        RECT  20.730 3.510 20.920 3.770 ;
        RECT  20.920 3.520 21.350 3.760 ;
        RECT  20.530 0.860 21.350 1.100 ;
        RECT  21.350 0.860 21.590 3.760 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.870 1.330 21.980 1.950 ;
        RECT  21.870 2.950 21.990 3.350 ;
        RECT  21.980 1.330 21.990 2.090 ;
        RECT  21.990 1.330 22.230 3.350 ;
        RECT  22.230 1.330 22.240 2.090 ;
        RECT  22.230 2.950 22.270 3.350 ;
        RECT  22.240 1.330 22.270 1.950 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.780 2.090 ;
        RECT  1.780 1.840 2.310 2.080 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.510 2.090 ;
        RECT  3.510 1.520 3.760 2.090 ;
        RECT  3.760 1.520 3.930 1.930 ;
        RECT  3.930 1.520 4.180 1.920 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.700 2.070 0.860 2.470 ;
        RECT  0.860 2.070 1.110 2.650 ;
        RECT  1.110 2.390 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.900 5.440 ;
        RECT  0.900 4.480 1.300 5.440 ;
        RECT  1.300 4.640 3.720 5.440 ;
        RECT  3.720 4.480 5.260 5.440 ;
        RECT  5.260 4.640 18.420 5.440 ;
        RECT  18.420 4.480 19.960 5.440 ;
        RECT  19.960 4.640 21.160 5.440 ;
        RECT  21.160 4.480 21.560 5.440 ;
        RECT  21.560 4.640 22.440 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.270 0.400 ;
        RECT  1.270 -0.400 2.320 0.560 ;
        RECT  2.320 -0.400 4.100 0.400 ;
        RECT  4.100 -0.400 4.500 0.560 ;
        RECT  4.500 -0.400 7.060 0.400 ;
        RECT  7.060 -0.400 7.460 0.560 ;
        RECT  7.460 -0.400 11.720 0.400 ;
        RECT  11.720 -0.400 11.960 1.050 ;
        RECT  11.960 -0.400 16.610 0.400 ;
        RECT  16.610 -0.400 17.010 0.910 ;
        RECT  17.010 -0.400 19.240 0.400 ;
        RECT  19.240 -0.400 19.250 0.750 ;
        RECT  19.250 -0.400 19.650 0.870 ;
        RECT  19.650 -0.400 19.660 0.750 ;
        RECT  19.660 -0.400 20.950 0.400 ;
        RECT  20.950 -0.400 21.350 0.560 ;
        RECT  21.350 -0.400 22.440 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  20.770 1.980 21.070 2.380 ;
        RECT  20.770 2.770 20.830 3.170 ;
        RECT  20.540 1.570 20.770 3.170 ;
        RECT  20.530 1.410 20.540 3.170 ;
        RECT  20.140 1.410 20.530 1.810 ;
        RECT  20.430 2.770 20.530 3.170 ;
        RECT  20.200 2.930 20.430 3.170 ;
        RECT  19.960 2.930 20.200 4.170 ;
        RECT  18.150 3.930 19.960 4.170 ;
        RECT  19.440 1.150 19.680 3.490 ;
        RECT  18.960 1.150 19.440 1.390 ;
        RECT  18.770 3.250 19.440 3.490 ;
        RECT  18.920 1.670 19.160 2.400 ;
        RECT  18.720 1.070 18.960 1.390 ;
        RECT  18.070 1.670 18.920 1.910 ;
        RECT  18.370 3.250 18.770 3.650 ;
        RECT  18.230 1.070 18.720 1.310 ;
        RECT  18.120 2.430 18.520 2.960 ;
        RECT  17.630 3.410 18.370 3.650 ;
        RECT  17.990 0.910 18.230 1.310 ;
        RECT  17.910 3.930 18.150 4.360 ;
        RECT  17.110 2.720 18.120 2.960 ;
        RECT  17.710 1.640 18.070 1.910 ;
        RECT  5.770 4.120 17.910 4.360 ;
        RECT  17.470 1.150 17.710 2.440 ;
        RECT  17.390 3.410 17.630 3.840 ;
        RECT  16.050 1.150 17.470 1.390 ;
        RECT  16.590 2.200 17.470 2.440 ;
        RECT  16.710 3.600 17.390 3.840 ;
        RECT  15.960 1.670 17.190 1.910 ;
        RECT  16.870 2.720 17.110 3.320 ;
        RECT  16.430 3.080 16.870 3.320 ;
        RECT  16.350 2.200 16.590 2.800 ;
        RECT  16.190 3.080 16.430 3.680 ;
        RECT  16.190 2.560 16.350 2.800 ;
        RECT  16.080 3.440 16.190 3.680 ;
        RECT  15.840 3.440 16.080 3.840 ;
        RECT  15.810 0.680 16.050 1.390 ;
        RECT  15.910 1.670 15.960 2.130 ;
        RECT  15.720 1.670 15.910 3.160 ;
        RECT  6.570 3.600 15.840 3.840 ;
        RECT  12.480 0.680 15.810 0.920 ;
        RECT  15.670 1.890 15.720 3.160 ;
        RECT  15.010 2.920 15.670 3.160 ;
        RECT  15.390 1.200 15.440 1.600 ;
        RECT  15.200 1.200 15.390 2.640 ;
        RECT  15.150 1.210 15.200 2.640 ;
        RECT  13.640 1.210 15.150 1.450 ;
        RECT  13.850 2.400 15.150 2.640 ;
        RECT  14.770 2.920 15.010 3.320 ;
        RECT  14.630 1.720 14.870 2.120 ;
        RECT  9.080 3.080 14.770 3.320 ;
        RECT  13.240 1.720 14.630 1.960 ;
        RECT  13.610 2.400 13.850 2.800 ;
        RECT  11.410 2.560 13.610 2.800 ;
        RECT  13.000 1.200 13.240 1.960 ;
        RECT  12.760 1.200 13.000 1.440 ;
        RECT  10.920 1.850 12.630 2.250 ;
        RECT  12.240 0.680 12.480 1.570 ;
        RECT  11.440 1.330 12.240 1.570 ;
        RECT  11.200 0.670 11.440 1.570 ;
        RECT  7.980 0.670 11.200 0.910 ;
        RECT  10.680 1.190 10.920 2.800 ;
        RECT  10.110 1.190 10.680 1.430 ;
        RECT  9.760 2.560 10.680 2.800 ;
        RECT  9.360 2.230 9.760 2.800 ;
        RECT  8.840 1.200 9.080 3.320 ;
        RECT  8.650 1.200 8.840 1.440 ;
        RECT  7.910 2.930 8.840 3.320 ;
        RECT  8.160 1.710 8.560 2.110 ;
        RECT  6.180 1.710 8.160 1.950 ;
        RECT  7.740 0.670 7.980 1.110 ;
        RECT  7.090 2.930 7.910 3.170 ;
        RECT  6.700 0.870 7.740 1.110 ;
        RECT  6.850 2.230 7.090 3.170 ;
        RECT  6.690 2.230 6.850 2.630 ;
        RECT  6.460 0.670 6.700 1.110 ;
        RECT  6.330 3.410 6.570 3.840 ;
        RECT  6.210 0.670 6.460 0.910 ;
        RECT  5.470 3.410 6.330 3.650 ;
        RECT  6.110 1.190 6.180 1.950 ;
        RECT  5.990 1.190 6.110 2.710 ;
        RECT  5.870 1.190 5.990 3.130 ;
        RECT  5.750 2.470 5.870 3.130 ;
        RECT  5.530 3.940 5.770 4.360 ;
        RECT  5.470 1.500 5.580 1.740 ;
        RECT  2.250 3.940 5.530 4.180 ;
        RECT  5.230 1.500 5.470 3.650 ;
        RECT  3.420 0.940 5.380 1.180 ;
        RECT  5.180 1.500 5.230 1.740 ;
        RECT  0.490 3.410 5.230 3.650 ;
        RECT  4.670 2.140 4.910 2.610 ;
        RECT  2.910 2.890 4.790 3.130 ;
        RECT  2.850 2.370 4.670 2.610 ;
        RECT  3.180 0.790 3.420 1.180 ;
        RECT  2.760 0.790 3.180 1.030 ;
        RECT  2.610 1.310 2.850 2.610 ;
        RECT  2.110 1.310 2.610 1.550 ;
        RECT  2.570 2.370 2.610 2.610 ;
        RECT  2.330 2.370 2.570 3.070 ;
        RECT  2.170 2.830 2.330 3.070 ;
        RECT  1.710 1.150 2.110 1.550 ;
        RECT  0.410 1.150 0.570 1.550 ;
        RECT  0.410 2.750 0.490 3.650 ;
        RECT  0.250 1.150 0.410 3.650 ;
        RECT  0.170 1.150 0.250 3.250 ;
    END
END JKFFSRXL

MACRO JKFFSRX4
    CLASS CORE ;
    FOREIGN JKFFSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFSRXL ;
    SIZE 25.080 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.370 2.250 7.830 2.660 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.440 1.270 9.550 1.530 ;
        RECT  9.550 1.270 9.700 1.950 ;
        RECT  9.700 1.290 9.790 1.950 ;
        RECT  9.790 1.710 10.160 1.950 ;
        RECT  10.160 1.710 10.400 2.120 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.230 1.820 21.240 3.220 ;
        RECT  21.240 1.140 21.660 3.220 ;
        RECT  21.660 1.820 21.670 3.220 ;
        RECT  21.660 1.140 21.910 1.560 ;
        RECT  21.670 2.760 22.010 3.180 ;
        RECT  21.910 1.150 22.110 1.550 ;
        RECT  22.010 2.770 22.210 3.170 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  23.210 2.380 23.480 3.780 ;
        RECT  23.050 1.150 23.480 1.550 ;
        RECT  23.480 1.150 23.650 3.780 ;
        RECT  23.650 1.150 23.770 3.740 ;
        RECT  23.770 1.150 23.880 3.080 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.780 2.090 ;
        RECT  1.780 1.840 2.250 2.080 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.510 2.090 ;
        RECT  3.510 1.600 3.760 2.090 ;
        RECT  3.760 1.600 4.180 1.840 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.700 2.120 0.860 2.520 ;
        RECT  0.860 2.120 1.110 2.650 ;
        RECT  1.110 2.390 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.780 5.440 ;
        RECT  0.780 4.480 1.180 5.440 ;
        RECT  1.180 4.640 3.650 5.440 ;
        RECT  3.650 4.480 5.190 5.440 ;
        RECT  5.190 4.640 18.500 5.440 ;
        RECT  18.500 4.480 20.040 5.440 ;
        RECT  20.040 4.640 21.160 5.440 ;
        RECT  21.160 4.210 21.170 5.440 ;
        RECT  21.170 4.010 21.570 5.440 ;
        RECT  21.570 4.210 21.580 5.440 ;
        RECT  21.580 4.640 22.620 5.440 ;
        RECT  22.620 4.250 22.630 5.440 ;
        RECT  22.630 4.050 23.030 5.440 ;
        RECT  23.030 4.250 23.040 5.440 ;
        RECT  23.040 4.640 24.010 5.440 ;
        RECT  24.010 4.250 24.020 5.440 ;
        RECT  24.020 4.050 24.420 5.440 ;
        RECT  24.420 4.250 24.430 5.440 ;
        RECT  24.430 4.640 25.080 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.270 0.400 ;
        RECT  1.270 -0.400 2.320 0.560 ;
        RECT  2.320 -0.400 4.100 0.400 ;
        RECT  4.100 -0.400 4.500 0.560 ;
        RECT  4.500 -0.400 7.070 0.400 ;
        RECT  7.070 -0.400 7.470 0.560 ;
        RECT  7.470 -0.400 11.720 0.400 ;
        RECT  11.720 -0.400 11.960 1.050 ;
        RECT  11.960 -0.400 16.670 0.400 ;
        RECT  16.670 -0.400 16.680 0.840 ;
        RECT  16.680 -0.400 17.080 0.960 ;
        RECT  17.080 -0.400 17.090 0.840 ;
        RECT  17.090 -0.400 19.410 0.400 ;
        RECT  19.410 -0.400 19.420 0.810 ;
        RECT  19.420 -0.400 19.820 0.930 ;
        RECT  19.820 -0.400 19.830 0.810 ;
        RECT  19.830 -0.400 21.080 0.400 ;
        RECT  21.080 -0.400 21.090 0.670 ;
        RECT  21.090 -0.400 21.490 0.870 ;
        RECT  21.490 -0.400 21.500 0.670 ;
        RECT  21.500 -0.400 22.370 0.400 ;
        RECT  22.370 -0.400 22.380 0.670 ;
        RECT  22.380 -0.400 22.780 0.870 ;
        RECT  22.780 -0.400 22.790 0.670 ;
        RECT  22.790 -0.400 23.660 0.400 ;
        RECT  23.660 -0.400 23.670 0.670 ;
        RECT  23.670 -0.400 24.070 0.870 ;
        RECT  24.070 -0.400 24.080 0.670 ;
        RECT  24.080 -0.400 25.080 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  22.730 1.850 23.240 2.090 ;
        RECT  22.490 1.850 22.730 3.730 ;
        RECT  20.770 3.490 22.490 3.730 ;
        RECT  20.640 2.770 20.770 3.730 ;
        RECT  20.610 1.080 20.640 3.730 ;
        RECT  20.400 1.080 20.610 4.180 ;
        RECT  20.240 1.080 20.400 1.480 ;
        RECT  20.370 2.770 20.400 4.180 ;
        RECT  18.220 3.940 20.370 4.180 ;
        RECT  19.550 1.210 19.790 3.660 ;
        RECT  18.390 1.210 19.550 1.450 ;
        RECT  17.700 3.420 19.550 3.660 ;
        RECT  19.030 1.750 19.270 2.550 ;
        RECT  17.870 1.750 19.030 1.990 ;
        RECT  18.310 2.390 18.550 3.140 ;
        RECT  18.150 0.950 18.390 1.450 ;
        RECT  17.180 2.900 18.310 3.140 ;
        RECT  17.980 3.940 18.220 4.360 ;
        RECT  6.050 4.120 17.980 4.360 ;
        RECT  17.630 1.240 17.870 2.590 ;
        RECT  17.460 3.420 17.700 3.840 ;
        RECT  16.120 1.240 17.630 1.480 ;
        RECT  16.660 2.350 17.630 2.590 ;
        RECT  16.860 3.600 17.460 3.840 ;
        RECT  16.060 1.830 17.350 2.070 ;
        RECT  16.940 2.900 17.180 3.320 ;
        RECT  16.580 3.080 16.940 3.320 ;
        RECT  16.420 2.350 16.660 2.750 ;
        RECT  16.340 3.080 16.580 3.530 ;
        RECT  15.930 3.290 16.340 3.530 ;
        RECT  15.880 0.680 16.120 1.480 ;
        RECT  15.820 1.830 16.060 3.010 ;
        RECT  15.690 3.290 15.930 3.840 ;
        RECT  12.480 0.680 15.880 0.920 ;
        RECT  15.010 2.770 15.820 3.010 ;
        RECT  6.570 3.600 15.690 3.840 ;
        RECT  15.270 1.200 15.510 2.490 ;
        RECT  13.790 1.200 15.270 1.440 ;
        RECT  13.930 2.250 15.270 2.490 ;
        RECT  14.770 2.770 15.010 3.320 ;
        RECT  13.510 1.720 14.990 1.960 ;
        RECT  9.080 3.080 14.770 3.320 ;
        RECT  13.690 2.250 13.930 2.800 ;
        RECT  11.230 2.560 13.690 2.800 ;
        RECT  13.270 1.200 13.510 1.960 ;
        RECT  12.760 1.200 13.270 1.440 ;
        RECT  10.920 1.880 12.990 2.280 ;
        RECT  12.240 0.680 12.480 1.580 ;
        RECT  11.440 1.340 12.240 1.580 ;
        RECT  11.200 0.670 11.440 1.580 ;
        RECT  7.980 0.670 11.200 0.910 ;
        RECT  10.680 1.190 10.920 2.800 ;
        RECT  10.110 1.190 10.680 1.430 ;
        RECT  9.760 2.560 10.680 2.800 ;
        RECT  9.360 2.250 9.760 2.800 ;
        RECT  8.840 1.200 9.080 3.320 ;
        RECT  8.650 1.200 8.840 1.440 ;
        RECT  7.910 2.930 8.840 3.320 ;
        RECT  8.160 1.710 8.560 2.110 ;
        RECT  6.260 1.710 8.160 1.950 ;
        RECT  7.740 0.670 7.980 1.110 ;
        RECT  7.090 2.930 7.910 3.170 ;
        RECT  6.780 0.870 7.740 1.110 ;
        RECT  6.850 2.230 7.090 3.170 ;
        RECT  6.690 2.230 6.850 2.630 ;
        RECT  6.540 0.670 6.780 1.110 ;
        RECT  6.330 3.410 6.570 3.840 ;
        RECT  6.210 0.670 6.540 0.910 ;
        RECT  5.390 3.410 6.330 3.650 ;
        RECT  6.020 1.150 6.260 3.080 ;
        RECT  5.810 3.940 6.050 4.360 ;
        RECT  5.860 1.150 6.020 1.550 ;
        RECT  5.670 2.840 6.020 3.080 ;
        RECT  2.130 3.940 5.810 4.180 ;
        RECT  5.390 1.500 5.580 1.740 ;
        RECT  5.150 1.500 5.390 3.650 ;
        RECT  3.310 0.940 5.380 1.180 ;
        RECT  0.490 3.410 5.150 3.650 ;
        RECT  4.470 2.320 4.870 2.610 ;
        RECT  2.790 2.880 4.730 3.120 ;
        RECT  2.780 2.370 4.470 2.610 ;
        RECT  3.070 0.790 3.310 1.180 ;
        RECT  2.760 0.790 3.070 1.030 ;
        RECT  2.540 1.310 2.780 2.610 ;
        RECT  2.110 1.310 2.540 1.550 ;
        RECT  2.450 2.370 2.540 2.610 ;
        RECT  2.210 2.370 2.450 3.070 ;
        RECT  2.050 2.830 2.210 3.070 ;
        RECT  1.710 1.150 2.110 1.550 ;
        RECT  0.410 1.150 0.570 1.550 ;
        RECT  0.410 2.850 0.490 3.650 ;
        RECT  0.250 1.150 0.410 3.650 ;
        RECT  0.170 1.150 0.250 3.250 ;
    END
END JKFFSRX4

MACRO JKFFSRX2
    CLASS CORE ;
    FOREIGN JKFFSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFSRXL ;
    SIZE 23.100 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.370 2.250 7.830 2.660 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.440 1.270 9.550 1.530 ;
        RECT  9.550 1.270 9.700 1.950 ;
        RECT  9.700 1.290 9.790 1.950 ;
        RECT  9.790 1.710 10.160 1.950 ;
        RECT  10.160 1.710 10.400 2.120 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.060 2.920 21.120 3.320 ;
        RECT  20.960 0.920 21.120 1.320 ;
        RECT  21.120 0.920 21.360 3.320 ;
        RECT  21.360 2.920 21.460 3.320 ;
        RECT  21.360 1.830 21.580 2.090 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.980 1.270 22.000 1.530 ;
        RECT  22.000 1.260 22.400 1.530 ;
        RECT  22.500 2.980 22.680 3.960 ;
        RECT  22.400 1.040 22.680 1.530 ;
        RECT  22.680 1.040 22.800 3.960 ;
        RECT  22.800 1.290 22.900 3.960 ;
        RECT  22.900 1.290 22.920 3.230 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.780 2.090 ;
        RECT  1.780 1.840 2.250 2.080 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.510 2.090 ;
        RECT  3.510 1.600 3.760 2.090 ;
        RECT  3.760 1.600 4.180 1.840 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.700 2.120 0.860 2.520 ;
        RECT  0.860 2.120 1.110 2.650 ;
        RECT  1.110 2.390 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.780 5.440 ;
        RECT  0.780 4.480 1.180 5.440 ;
        RECT  1.180 4.640 3.650 5.440 ;
        RECT  3.650 4.480 5.190 5.440 ;
        RECT  5.190 4.640 18.470 5.440 ;
        RECT  18.470 4.480 20.010 5.440 ;
        RECT  20.010 4.640 21.770 5.440 ;
        RECT  21.770 4.320 21.780 5.440 ;
        RECT  21.780 4.120 22.180 5.440 ;
        RECT  22.180 4.320 22.190 5.440 ;
        RECT  22.190 4.640 23.100 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.270 0.400 ;
        RECT  1.270 -0.400 2.320 0.560 ;
        RECT  2.320 -0.400 4.100 0.400 ;
        RECT  4.100 -0.400 4.500 0.560 ;
        RECT  4.500 -0.400 7.070 0.400 ;
        RECT  7.070 -0.400 7.470 0.560 ;
        RECT  7.470 -0.400 11.720 0.400 ;
        RECT  11.720 -0.400 11.960 1.050 ;
        RECT  11.960 -0.400 16.640 0.400 ;
        RECT  16.640 -0.400 16.650 0.840 ;
        RECT  16.650 -0.400 17.050 0.960 ;
        RECT  17.050 -0.400 17.060 0.840 ;
        RECT  17.060 -0.400 19.380 0.400 ;
        RECT  19.380 -0.400 19.390 0.810 ;
        RECT  19.390 -0.400 19.790 0.930 ;
        RECT  19.790 -0.400 19.800 0.810 ;
        RECT  19.800 -0.400 21.670 0.400 ;
        RECT  21.670 -0.400 21.680 0.790 ;
        RECT  21.680 -0.400 22.080 0.990 ;
        RECT  22.080 -0.400 22.090 0.790 ;
        RECT  22.090 -0.400 23.100 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  22.000 2.260 22.400 2.660 ;
        RECT  21.980 2.420 22.000 2.660 ;
        RECT  21.740 2.420 21.980 3.840 ;
        RECT  20.800 3.600 21.740 3.840 ;
        RECT  20.610 3.600 20.800 4.180 ;
        RECT  20.370 1.080 20.610 4.180 ;
        RECT  20.210 1.080 20.370 1.480 ;
        RECT  18.190 3.940 20.370 4.180 ;
        RECT  19.520 1.210 19.760 3.660 ;
        RECT  18.360 1.210 19.520 1.450 ;
        RECT  17.670 3.420 19.520 3.660 ;
        RECT  19.000 1.750 19.240 2.550 ;
        RECT  17.840 1.750 19.000 1.990 ;
        RECT  18.280 2.390 18.520 3.140 ;
        RECT  18.120 0.950 18.360 1.450 ;
        RECT  17.150 2.900 18.280 3.140 ;
        RECT  17.950 3.940 18.190 4.360 ;
        RECT  6.050 4.120 17.950 4.360 ;
        RECT  17.600 1.240 17.840 2.590 ;
        RECT  17.430 3.420 17.670 3.840 ;
        RECT  16.090 1.240 17.600 1.480 ;
        RECT  16.630 2.350 17.600 2.590 ;
        RECT  16.830 3.600 17.430 3.840 ;
        RECT  16.030 1.830 17.320 2.070 ;
        RECT  16.910 2.900 17.150 3.320 ;
        RECT  16.550 3.080 16.910 3.320 ;
        RECT  16.390 2.350 16.630 2.750 ;
        RECT  16.310 3.080 16.550 3.530 ;
        RECT  15.980 3.290 16.310 3.530 ;
        RECT  15.850 0.680 16.090 1.480 ;
        RECT  15.790 1.830 16.030 3.010 ;
        RECT  15.740 3.290 15.980 3.840 ;
        RECT  12.480 0.680 15.850 0.920 ;
        RECT  15.010 2.770 15.790 3.010 ;
        RECT  6.570 3.600 15.740 3.840 ;
        RECT  15.270 1.200 15.510 2.490 ;
        RECT  13.720 1.200 15.270 1.440 ;
        RECT  13.930 2.250 15.270 2.490 ;
        RECT  14.770 2.770 15.010 3.320 ;
        RECT  13.440 1.720 14.990 1.960 ;
        RECT  9.080 3.080 14.770 3.320 ;
        RECT  13.690 2.250 13.930 2.800 ;
        RECT  11.230 2.560 13.690 2.800 ;
        RECT  13.200 1.200 13.440 1.960 ;
        RECT  12.760 1.200 13.200 1.440 ;
        RECT  10.920 1.880 12.920 2.280 ;
        RECT  12.240 0.680 12.480 1.580 ;
        RECT  11.440 1.340 12.240 1.580 ;
        RECT  11.200 0.670 11.440 1.580 ;
        RECT  7.980 0.670 11.200 0.910 ;
        RECT  10.680 1.190 10.920 2.800 ;
        RECT  10.110 1.190 10.680 1.430 ;
        RECT  9.760 2.560 10.680 2.800 ;
        RECT  9.360 2.250 9.760 2.800 ;
        RECT  8.840 1.190 9.080 3.320 ;
        RECT  8.650 1.190 8.840 1.430 ;
        RECT  7.910 2.930 8.840 3.320 ;
        RECT  8.160 1.710 8.560 2.110 ;
        RECT  6.260 1.710 8.160 1.950 ;
        RECT  7.740 0.670 7.980 1.110 ;
        RECT  7.090 2.930 7.910 3.170 ;
        RECT  6.780 0.870 7.740 1.110 ;
        RECT  6.850 2.230 7.090 3.170 ;
        RECT  6.690 2.230 6.850 2.630 ;
        RECT  6.540 0.670 6.780 1.110 ;
        RECT  6.330 3.410 6.570 3.840 ;
        RECT  6.210 0.670 6.540 0.910 ;
        RECT  5.390 3.410 6.330 3.650 ;
        RECT  6.020 1.150 6.260 3.080 ;
        RECT  5.810 3.940 6.050 4.360 ;
        RECT  5.860 1.150 6.020 1.550 ;
        RECT  5.670 2.840 6.020 3.080 ;
        RECT  2.130 3.940 5.810 4.180 ;
        RECT  5.390 1.500 5.580 1.740 ;
        RECT  5.150 1.500 5.390 3.650 ;
        RECT  3.310 0.940 5.380 1.180 ;
        RECT  0.490 3.410 5.150 3.650 ;
        RECT  4.470 2.320 4.870 2.610 ;
        RECT  2.790 2.880 4.730 3.120 ;
        RECT  2.780 2.370 4.470 2.610 ;
        RECT  3.070 0.790 3.310 1.180 ;
        RECT  2.760 0.790 3.070 1.030 ;
        RECT  2.540 1.310 2.780 2.610 ;
        RECT  2.110 1.310 2.540 1.550 ;
        RECT  2.450 2.370 2.540 2.610 ;
        RECT  2.210 2.370 2.450 3.070 ;
        RECT  2.050 2.830 2.210 3.070 ;
        RECT  1.710 1.150 2.110 1.550 ;
        RECT  0.410 1.150 0.570 1.550 ;
        RECT  0.410 2.850 0.490 3.650 ;
        RECT  0.250 1.150 0.410 3.650 ;
        RECT  0.170 1.150 0.250 3.250 ;
    END
END JKFFSRX2

MACRO JKFFSRX1
    CLASS CORE ;
    FOREIGN JKFFSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFSRXL ;
    SIZE 22.440 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.370 2.250 7.830 2.660 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.440 1.270 9.550 1.530 ;
        RECT  9.550 1.270 9.700 1.950 ;
        RECT  9.700 1.290 9.790 1.950 ;
        RECT  9.790 1.710 10.160 1.950 ;
        RECT  10.160 1.710 10.400 2.120 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  20.070 0.670 20.470 1.100 ;
        RECT  20.490 3.520 20.660 4.340 ;
        RECT  20.660 3.510 20.730 4.340 ;
        RECT  20.730 3.510 20.920 3.770 ;
        RECT  20.920 3.520 21.350 3.760 ;
        RECT  20.470 0.860 21.350 1.100 ;
        RECT  21.350 0.860 21.590 3.760 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.870 1.340 21.980 1.960 ;
        RECT  21.870 2.920 21.990 3.320 ;
        RECT  21.980 1.340 21.990 2.090 ;
        RECT  21.990 1.340 22.230 3.320 ;
        RECT  22.230 1.340 22.240 2.090 ;
        RECT  22.230 2.920 22.270 3.320 ;
        RECT  22.240 1.340 22.270 1.960 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.780 2.090 ;
        RECT  1.780 1.840 2.250 2.080 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.510 2.090 ;
        RECT  3.510 1.600 3.760 2.090 ;
        RECT  3.760 1.600 4.180 1.840 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.700 2.120 0.860 2.520 ;
        RECT  0.860 2.120 1.110 2.650 ;
        RECT  1.110 2.390 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.780 5.440 ;
        RECT  0.780 4.480 1.180 5.440 ;
        RECT  1.180 4.640 3.660 5.440 ;
        RECT  3.660 4.480 5.200 5.440 ;
        RECT  5.200 4.640 18.420 5.440 ;
        RECT  18.420 4.480 19.960 5.440 ;
        RECT  19.960 4.640 21.140 5.440 ;
        RECT  21.140 4.480 21.540 5.440 ;
        RECT  21.540 4.640 22.440 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.270 0.400 ;
        RECT  1.270 -0.400 2.320 0.560 ;
        RECT  2.320 -0.400 4.100 0.400 ;
        RECT  4.100 -0.400 4.500 0.560 ;
        RECT  4.500 -0.400 7.060 0.400 ;
        RECT  7.060 -0.400 7.460 0.560 ;
        RECT  7.460 -0.400 11.720 0.400 ;
        RECT  11.720 -0.400 11.960 1.050 ;
        RECT  11.960 -0.400 16.600 0.400 ;
        RECT  16.600 -0.400 16.610 0.750 ;
        RECT  16.610 -0.400 17.010 0.870 ;
        RECT  17.010 -0.400 17.020 0.750 ;
        RECT  17.020 -0.400 19.240 0.400 ;
        RECT  19.240 -0.400 19.250 0.750 ;
        RECT  19.250 -0.400 19.650 0.870 ;
        RECT  19.650 -0.400 19.660 0.750 ;
        RECT  19.660 -0.400 21.010 0.400 ;
        RECT  21.010 -0.400 21.410 0.560 ;
        RECT  21.410 -0.400 22.440 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  20.770 1.980 21.070 2.380 ;
        RECT  20.530 1.570 20.770 3.170 ;
        RECT  20.480 1.570 20.530 1.810 ;
        RECT  20.370 2.770 20.530 3.170 ;
        RECT  20.080 1.410 20.480 1.810 ;
        RECT  20.210 2.930 20.370 3.170 ;
        RECT  19.970 2.930 20.210 4.170 ;
        RECT  18.150 3.930 19.970 4.170 ;
        RECT  19.440 1.150 19.680 3.490 ;
        RECT  18.960 1.150 19.440 1.390 ;
        RECT  18.770 3.250 19.440 3.490 ;
        RECT  18.920 1.670 19.160 2.400 ;
        RECT  18.720 1.070 18.960 1.390 ;
        RECT  18.070 1.670 18.920 1.910 ;
        RECT  18.370 3.250 18.770 3.650 ;
        RECT  18.230 1.070 18.720 1.310 ;
        RECT  18.120 2.430 18.520 2.960 ;
        RECT  17.630 3.410 18.370 3.650 ;
        RECT  17.990 0.910 18.230 1.310 ;
        RECT  17.910 3.930 18.150 4.360 ;
        RECT  17.110 2.720 18.120 2.960 ;
        RECT  17.710 1.600 18.070 1.910 ;
        RECT  6.050 4.120 17.910 4.360 ;
        RECT  17.470 1.150 17.710 2.440 ;
        RECT  17.390 3.410 17.630 3.840 ;
        RECT  16.050 1.150 17.470 1.390 ;
        RECT  16.590 2.200 17.470 2.440 ;
        RECT  16.710 3.600 17.390 3.840 ;
        RECT  15.960 1.670 17.190 1.910 ;
        RECT  16.870 2.720 17.110 3.320 ;
        RECT  16.430 3.080 16.870 3.320 ;
        RECT  16.350 2.200 16.590 2.800 ;
        RECT  16.190 3.080 16.430 3.680 ;
        RECT  16.190 2.560 16.350 2.800 ;
        RECT  16.080 3.440 16.190 3.680 ;
        RECT  15.840 3.440 16.080 3.840 ;
        RECT  15.810 0.680 16.050 1.390 ;
        RECT  15.910 1.670 15.960 2.130 ;
        RECT  15.720 1.670 15.910 3.160 ;
        RECT  6.570 3.600 15.840 3.840 ;
        RECT  12.480 0.680 15.810 0.920 ;
        RECT  15.670 1.890 15.720 3.160 ;
        RECT  15.010 2.920 15.670 3.160 ;
        RECT  15.390 1.200 15.440 1.600 ;
        RECT  15.150 1.200 15.390 2.640 ;
        RECT  13.520 1.200 15.150 1.440 ;
        RECT  13.850 2.400 15.150 2.640 ;
        RECT  14.770 2.920 15.010 3.320 ;
        RECT  14.630 1.720 14.870 2.120 ;
        RECT  9.080 3.080 14.770 3.320 ;
        RECT  13.220 1.720 14.630 1.960 ;
        RECT  13.610 2.400 13.850 2.800 ;
        RECT  11.470 2.560 13.610 2.800 ;
        RECT  12.980 1.200 13.220 1.960 ;
        RECT  12.760 1.200 12.980 1.440 ;
        RECT  10.920 1.850 12.630 2.250 ;
        RECT  12.240 0.680 12.480 1.570 ;
        RECT  11.440 1.330 12.240 1.570 ;
        RECT  11.200 0.670 11.440 1.570 ;
        RECT  7.980 0.670 11.200 0.910 ;
        RECT  10.680 1.190 10.920 2.800 ;
        RECT  10.110 1.190 10.680 1.430 ;
        RECT  9.760 2.560 10.680 2.800 ;
        RECT  9.360 2.250 9.760 2.800 ;
        RECT  8.840 1.190 9.080 3.320 ;
        RECT  8.650 1.190 8.840 1.430 ;
        RECT  7.910 2.920 8.840 3.320 ;
        RECT  8.160 1.710 8.560 2.110 ;
        RECT  6.180 1.710 8.160 1.950 ;
        RECT  7.740 0.670 7.980 1.110 ;
        RECT  7.090 2.920 7.910 3.160 ;
        RECT  6.730 0.870 7.740 1.110 ;
        RECT  6.850 2.230 7.090 3.160 ;
        RECT  6.690 2.230 6.850 2.630 ;
        RECT  6.490 0.670 6.730 1.110 ;
        RECT  6.330 3.410 6.570 3.840 ;
        RECT  6.210 0.670 6.490 0.910 ;
        RECT  5.390 3.410 6.330 3.650 ;
        RECT  5.940 1.150 6.180 3.080 ;
        RECT  5.810 3.940 6.050 4.360 ;
        RECT  5.670 2.840 5.940 3.080 ;
        RECT  2.130 3.940 5.810 4.180 ;
        RECT  5.390 1.500 5.580 1.740 ;
        RECT  5.150 1.500 5.390 3.650 ;
        RECT  3.310 0.940 5.380 1.180 ;
        RECT  0.490 3.410 5.150 3.650 ;
        RECT  4.470 2.320 4.870 2.610 ;
        RECT  2.790 2.880 4.730 3.120 ;
        RECT  2.780 2.370 4.470 2.610 ;
        RECT  3.070 0.790 3.310 1.180 ;
        RECT  2.760 0.790 3.070 1.030 ;
        RECT  2.540 1.310 2.780 2.610 ;
        RECT  2.110 1.310 2.540 1.550 ;
        RECT  2.450 2.370 2.540 2.610 ;
        RECT  2.210 2.370 2.450 3.070 ;
        RECT  2.050 2.830 2.210 3.070 ;
        RECT  1.710 1.150 2.110 1.550 ;
        RECT  0.410 1.150 0.570 1.550 ;
        RECT  0.410 2.850 0.490 3.650 ;
        RECT  0.250 1.150 0.410 3.650 ;
        RECT  0.170 1.150 0.250 3.250 ;
    END
END JKFFSRX1

MACRO JKFFSXL
    CLASS CORE ;
    FOREIGN JKFFSXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.820 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.780 1.650 8.050 1.890 ;
        RECT  8.050 0.670 8.290 1.890 ;
        RECT  8.290 0.670 12.620 0.910 ;
        RECT  12.620 0.670 12.860 1.100 ;
        RECT  12.860 0.860 13.820 1.100 ;
        RECT  13.820 0.670 14.220 1.100 ;
        RECT  14.220 0.710 14.320 0.970 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.600 2.970 15.880 3.410 ;
        RECT  15.580 1.390 15.880 1.790 ;
        RECT  15.880 1.390 15.980 3.410 ;
        RECT  15.980 1.470 16.000 3.410 ;
        RECT  16.000 1.470 16.120 3.210 ;
        RECT  16.120 2.950 16.300 3.210 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.250 2.950 17.370 3.350 ;
        RECT  17.360 2.390 17.370 2.650 ;
        RECT  17.250 1.380 17.370 1.950 ;
        RECT  17.370 1.380 17.610 3.350 ;
        RECT  17.610 2.390 17.620 2.650 ;
        RECT  17.610 2.950 17.650 3.350 ;
        RECT  17.610 1.380 17.650 1.950 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.780 2.090 ;
        RECT  1.780 1.850 2.310 2.090 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.070 1.690 4.540 2.100 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.710 2.070 0.860 2.470 ;
        RECT  0.860 2.070 1.110 2.650 ;
        RECT  1.110 2.390 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.880 5.440 ;
        RECT  0.880 4.480 1.280 5.440 ;
        RECT  1.280 4.640 3.980 5.440 ;
        RECT  3.980 4.480 4.380 5.440 ;
        RECT  4.380 4.640 6.940 5.440 ;
        RECT  6.940 4.480 7.920 5.440 ;
        RECT  7.920 4.640 14.210 5.440 ;
        RECT  14.210 4.480 15.190 5.440 ;
        RECT  15.190 4.640 16.420 5.440 ;
        RECT  16.420 4.480 16.820 5.440 ;
        RECT  16.820 4.640 17.820 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 2.370 0.400 ;
        RECT  2.370 -0.400 2.770 0.560 ;
        RECT  2.770 -0.400 4.440 0.400 ;
        RECT  4.440 -0.400 4.840 0.560 ;
        RECT  4.840 -0.400 7.360 0.400 ;
        RECT  7.360 -0.400 7.370 1.160 ;
        RECT  7.370 -0.400 7.770 1.360 ;
        RECT  7.770 -0.400 7.780 1.160 ;
        RECT  7.780 -0.400 13.140 0.400 ;
        RECT  13.140 -0.400 13.540 0.560 ;
        RECT  13.540 -0.400 16.470 0.400 ;
        RECT  16.470 -0.400 16.870 0.560 ;
        RECT  16.870 -0.400 17.820 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.970 2.190 17.000 2.590 ;
        RECT  16.730 0.860 16.970 4.180 ;
        RECT  15.980 0.860 16.730 1.100 ;
        RECT  15.940 3.940 16.730 4.180 ;
        RECT  15.580 0.670 15.980 1.100 ;
        RECT  15.540 3.940 15.940 4.350 ;
        RECT  13.640 3.940 15.540 4.180 ;
        RECT  15.180 2.130 15.380 2.530 ;
        RECT  15.180 1.160 15.240 1.560 ;
        RECT  14.940 1.160 15.180 3.650 ;
        RECT  14.840 1.160 14.940 1.620 ;
        RECT  14.060 3.410 14.940 3.650 ;
        RECT  13.360 1.380 14.840 1.620 ;
        RECT  13.120 2.650 14.660 3.050 ;
        RECT  13.400 3.940 13.640 4.360 ;
        RECT  8.430 4.120 13.400 4.360 ;
        RECT  13.120 1.380 13.360 2.140 ;
        RECT  12.880 2.430 13.120 3.750 ;
        RECT  12.840 2.430 12.880 2.670 ;
        RECT  11.960 3.510 12.880 3.750 ;
        RECT  12.600 1.390 12.840 2.670 ;
        RECT  12.340 1.390 12.600 1.630 ;
        RECT  12.320 2.950 12.600 3.190 ;
        RECT  12.100 1.190 12.340 1.630 ;
        RECT  12.080 1.910 12.320 3.190 ;
        RECT  11.680 1.190 12.100 1.430 ;
        RECT  11.820 1.910 12.080 2.150 ;
        RECT  11.430 1.790 11.820 2.150 ;
        RECT  11.680 2.430 11.800 2.830 ;
        RECT  11.440 2.430 11.680 3.830 ;
        RECT  10.670 2.430 11.440 2.670 ;
        RECT  8.950 3.590 11.440 3.830 ;
        RECT  11.190 1.790 11.430 2.030 ;
        RECT  10.950 1.190 11.190 2.030 ;
        RECT  11.070 2.950 11.150 3.190 ;
        RECT  10.750 2.950 11.070 3.310 ;
        RECT  9.860 1.190 10.950 1.430 ;
        RECT  9.470 3.070 10.750 3.310 ;
        RECT  10.580 1.790 10.670 2.670 ;
        RECT  10.430 1.710 10.580 2.670 ;
        RECT  10.340 1.710 10.430 2.110 ;
        RECT  9.990 2.550 10.150 2.790 ;
        RECT  9.860 1.760 9.990 2.790 ;
        RECT  9.750 1.190 9.860 2.790 ;
        RECT  9.620 1.190 9.750 2.080 ;
        RECT  9.340 2.810 9.470 3.310 ;
        RECT  9.230 1.190 9.340 3.310 ;
        RECT  9.100 1.190 9.230 3.050 ;
        RECT  8.800 1.190 9.100 1.430 ;
        RECT  7.740 2.810 9.100 3.050 ;
        RECT  8.710 3.420 8.950 3.830 ;
        RECT  8.580 1.710 8.820 2.410 ;
        RECT  6.940 3.420 8.710 3.660 ;
        RECT  7.460 2.170 8.580 2.410 ;
        RECT  8.190 3.940 8.430 4.360 ;
        RECT  3.590 3.940 8.190 4.180 ;
        RECT  7.340 2.690 7.740 3.050 ;
        RECT  7.220 2.030 7.460 2.410 ;
        RECT  6.370 2.030 7.220 2.270 ;
        RECT  6.700 2.610 6.940 3.660 ;
        RECT  5.770 3.420 6.700 3.660 ;
        RECT  6.370 1.010 6.430 1.410 ;
        RECT  6.130 1.010 6.370 3.140 ;
        RECT  6.030 1.010 6.130 1.410 ;
        RECT  5.750 1.680 5.770 3.660 ;
        RECT  5.530 1.570 5.750 3.660 ;
        RECT  3.510 1.050 5.550 1.290 ;
        RECT  5.350 1.570 5.530 1.970 ;
        RECT  2.890 2.890 5.530 3.130 ;
        RECT  2.830 2.370 5.250 2.610 ;
        RECT  3.170 3.410 5.110 3.650 ;
        RECT  3.170 3.940 3.590 4.220 ;
        RECT  3.110 1.000 3.510 1.400 ;
        RECT  2.610 3.980 3.170 4.220 ;
        RECT  2.650 2.890 2.890 3.670 ;
        RECT  2.590 1.230 2.830 2.610 ;
        RECT  0.490 3.430 2.650 3.670 ;
        RECT  1.710 1.230 2.590 1.470 ;
        RECT  2.370 2.370 2.590 2.610 ;
        RECT  2.130 2.370 2.370 3.150 ;
        RECT  0.410 1.220 0.570 1.620 ;
        RECT  0.410 2.750 0.490 3.670 ;
        RECT  0.250 1.220 0.410 3.670 ;
        RECT  0.170 1.220 0.250 3.190 ;
    END
END JKFFSXL

MACRO JKFFSX4
    CLASS CORE ;
    FOREIGN JKFFSX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFSXL ;
    SIZE 21.780 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.720 1.560 8.020 1.960 ;
        RECT  8.020 0.680 8.260 1.960 ;
        RECT  8.260 0.680 10.280 0.920 ;
        RECT  10.280 0.680 10.520 1.100 ;
        RECT  10.520 0.860 11.480 1.100 ;
        RECT  11.480 0.680 11.720 1.100 ;
        RECT  11.720 0.680 13.580 0.920 ;
        RECT  13.580 0.680 13.820 1.100 ;
        RECT  13.820 0.860 15.380 1.100 ;
        RECT  15.380 0.710 15.640 1.100 ;
        RECT  15.640 0.860 16.420 1.100 ;
        RECT  16.420 0.860 16.660 2.400 ;
        RECT  16.660 2.000 16.820 2.400 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.590 1.820 18.760 3.220 ;
        RECT  18.760 1.530 18.770 3.260 ;
        RECT  18.770 1.330 19.170 3.260 ;
        RECT  19.170 1.530 19.180 3.260 ;
        RECT  19.180 2.850 19.240 3.250 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  19.910 1.820 20.100 3.220 ;
        RECT  20.100 1.530 20.110 3.220 ;
        RECT  20.110 1.330 20.380 3.220 ;
        RECT  20.380 1.330 20.510 3.250 ;
        RECT  20.510 1.530 20.520 3.250 ;
        RECT  20.520 2.840 20.770 3.250 ;
        RECT  20.770 2.850 20.780 3.250 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.860 2.090 ;
        RECT  1.860 1.690 2.260 2.090 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.060 1.690 4.510 2.100 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.700 2.170 1.120 2.660 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.980 5.440 ;
        RECT  0.980 4.480 1.380 5.440 ;
        RECT  1.380 4.640 4.000 5.440 ;
        RECT  4.000 4.480 4.400 5.440 ;
        RECT  4.400 4.640 6.970 5.440 ;
        RECT  6.970 4.480 7.950 5.440 ;
        RECT  7.950 4.640 14.360 5.440 ;
        RECT  14.360 4.480 16.460 5.440 ;
        RECT  16.460 4.640 18.060 5.440 ;
        RECT  18.060 4.280 18.070 5.440 ;
        RECT  18.070 4.080 18.470 5.440 ;
        RECT  18.470 4.280 18.480 5.440 ;
        RECT  18.480 4.640 19.600 5.440 ;
        RECT  19.600 4.280 19.610 5.440 ;
        RECT  19.610 4.080 20.010 5.440 ;
        RECT  20.010 4.280 20.020 5.440 ;
        RECT  20.020 4.640 20.990 5.440 ;
        RECT  20.990 4.280 21.000 5.440 ;
        RECT  21.000 4.080 21.400 5.440 ;
        RECT  21.400 4.280 21.410 5.440 ;
        RECT  21.410 4.640 21.780 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.150 0.400 ;
        RECT  1.150 -0.400 1.230 0.560 ;
        RECT  1.230 -0.400 2.350 0.580 ;
        RECT  2.350 -0.400 2.720 0.560 ;
        RECT  2.720 -0.400 4.290 0.400 ;
        RECT  4.290 -0.400 4.690 0.560 ;
        RECT  4.690 -0.400 7.340 0.400 ;
        RECT  7.340 -0.400 7.740 1.320 ;
        RECT  7.740 -0.400 10.800 0.400 ;
        RECT  10.800 -0.400 11.200 0.560 ;
        RECT  11.200 -0.400 14.100 0.400 ;
        RECT  14.100 -0.400 14.500 0.560 ;
        RECT  14.500 -0.400 16.740 0.400 ;
        RECT  16.740 -0.400 17.140 0.560 ;
        RECT  17.140 -0.400 18.090 0.400 ;
        RECT  18.090 -0.400 18.100 0.850 ;
        RECT  18.100 -0.400 18.500 1.050 ;
        RECT  18.500 -0.400 18.510 0.850 ;
        RECT  18.510 -0.400 19.430 0.400 ;
        RECT  19.430 -0.400 19.440 0.850 ;
        RECT  19.440 -0.400 19.840 1.050 ;
        RECT  19.840 -0.400 19.850 0.850 ;
        RECT  19.850 -0.400 20.720 0.400 ;
        RECT  20.720 -0.400 20.730 0.850 ;
        RECT  20.730 -0.400 21.130 1.050 ;
        RECT  21.130 -0.400 21.140 0.850 ;
        RECT  21.140 -0.400 21.780 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  21.060 2.330 21.300 3.770 ;
        RECT  21.030 2.330 21.060 2.570 ;
        RECT  18.320 3.530 21.060 3.770 ;
        RECT  20.790 2.170 21.030 2.570 ;
        RECT  18.080 1.490 18.320 3.770 ;
        RECT  17.880 1.490 18.080 1.730 ;
        RECT  17.350 3.240 18.080 3.640 ;
        RECT  17.480 1.330 17.880 1.730 ;
        RECT  17.640 2.070 17.800 2.470 ;
        RECT  17.400 2.070 17.640 2.960 ;
        RECT  16.400 2.720 17.400 2.960 ;
        RECT  17.200 3.400 17.350 3.640 ;
        RECT  16.960 3.400 17.200 4.180 ;
        RECT  14.070 3.940 16.960 4.180 ;
        RECT  16.200 2.720 16.400 3.660 ;
        RECT  16.170 2.720 16.200 3.670 ;
        RECT  16.140 2.710 16.170 3.670 ;
        RECT  15.900 1.540 16.140 3.670 ;
        RECT  15.780 1.540 15.900 1.780 ;
        RECT  14.760 3.250 15.900 3.670 ;
        RECT  15.380 1.380 15.780 1.780 ;
        RECT  15.260 2.160 15.660 2.560 ;
        RECT  14.150 1.540 15.380 1.780 ;
        RECT  13.550 2.320 15.260 2.560 ;
        RECT  14.560 3.260 14.760 3.660 ;
        RECT  13.910 1.540 14.150 2.030 ;
        RECT  13.830 3.940 14.070 4.360 ;
        RECT  8.460 4.120 13.830 4.360 ;
        RECT  13.310 1.790 13.550 3.840 ;
        RECT  13.300 1.790 13.310 2.030 ;
        RECT  12.460 3.600 13.310 3.840 ;
        RECT  13.060 1.200 13.300 2.030 ;
        RECT  12.740 1.200 13.060 1.440 ;
        RECT  12.790 2.360 13.030 3.320 ;
        RECT  12.780 2.360 12.790 2.600 ;
        RECT  12.540 1.760 12.780 2.600 ;
        RECT  12.460 1.760 12.540 2.000 ;
        RECT  12.220 1.380 12.460 2.000 ;
        RECT  12.220 2.900 12.460 3.880 ;
        RECT  10.030 1.380 12.220 1.620 ;
        RECT  11.940 2.360 12.140 2.600 ;
        RECT  11.700 1.900 11.940 3.840 ;
        RECT  10.300 1.900 11.700 2.140 ;
        RECT  8.980 3.600 11.700 3.840 ;
        RECT  11.260 2.420 11.420 2.660 ;
        RECT  11.020 2.420 11.260 3.320 ;
        RECT  9.500 3.080 11.020 3.320 ;
        RECT  10.020 2.560 10.260 2.800 ;
        RECT  10.020 1.380 10.030 1.940 ;
        RECT  10.000 1.380 10.020 2.800 ;
        RECT  9.780 1.200 10.000 2.800 ;
        RECT  9.580 1.200 9.780 2.090 ;
        RECT  9.300 2.890 9.500 3.320 ;
        RECT  9.260 1.200 9.300 3.320 ;
        RECT  9.060 1.200 9.260 3.130 ;
        RECT  8.740 1.200 9.060 1.440 ;
        RECT  7.280 2.860 9.060 3.130 ;
        RECT  8.740 3.420 8.980 3.840 ;
        RECT  8.540 1.810 8.780 2.580 ;
        RECT  6.880 3.420 8.740 3.660 ;
        RECT  7.400 2.340 8.540 2.580 ;
        RECT  8.220 3.940 8.460 4.360 ;
        RECT  3.410 3.940 8.220 4.180 ;
        RECT  7.160 2.250 7.400 2.580 ;
        RECT  6.310 2.250 7.160 2.490 ;
        RECT  6.640 2.770 6.880 3.660 ;
        RECT  5.740 3.420 6.640 3.660 ;
        RECT  6.310 0.940 6.400 1.340 ;
        RECT  6.070 0.940 6.310 3.140 ;
        RECT  6.000 0.940 6.070 1.340 ;
        RECT  5.500 1.620 5.740 3.660 ;
        RECT  3.460 1.060 5.520 1.300 ;
        RECT  5.320 1.620 5.500 1.860 ;
        RECT  2.890 2.890 5.500 3.130 ;
        RECT  2.780 2.370 5.220 2.610 ;
        RECT  3.170 3.410 5.110 3.650 ;
        RECT  3.060 1.020 3.460 1.420 ;
        RECT  3.170 3.940 3.410 4.230 ;
        RECT  2.370 3.990 3.170 4.230 ;
        RECT  2.650 2.890 2.890 3.670 ;
        RECT  2.540 1.180 2.780 2.610 ;
        RECT  0.570 3.430 2.650 3.670 ;
        RECT  1.650 1.180 2.540 1.420 ;
        RECT  2.370 2.370 2.540 2.610 ;
        RECT  2.130 2.370 2.370 3.150 ;
        RECT  0.400 1.270 0.570 1.670 ;
        RECT  0.400 2.960 0.570 3.670 ;
        RECT  0.330 1.270 0.400 3.670 ;
        RECT  0.170 1.270 0.330 3.360 ;
        RECT  0.160 1.280 0.170 3.350 ;
    END
END JKFFSX4

MACRO JKFFSX2
    CLASS CORE ;
    FOREIGN JKFFSX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFSXL ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.780 1.650 8.050 1.890 ;
        RECT  8.050 0.670 8.290 1.890 ;
        RECT  8.290 0.670 12.620 0.910 ;
        RECT  12.620 0.670 12.860 1.100 ;
        RECT  12.860 0.860 13.980 1.100 ;
        RECT  13.980 0.670 14.300 1.100 ;
        RECT  14.300 0.670 14.320 0.970 ;
        RECT  14.320 0.670 15.330 0.910 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.290 2.850 16.610 3.250 ;
        RECT  16.630 1.540 16.640 2.100 ;
        RECT  16.610 2.660 16.680 3.250 ;
        RECT  16.640 1.360 16.680 2.100 ;
        RECT  16.680 1.360 16.690 3.250 ;
        RECT  16.690 1.360 16.710 3.200 ;
        RECT  16.710 1.360 16.920 3.090 ;
        RECT  16.920 1.360 17.040 2.100 ;
        RECT  17.040 1.540 17.050 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.320 1.520 17.560 3.260 ;
        RECT  17.560 2.860 17.850 3.260 ;
        RECT  17.560 1.520 17.880 1.760 ;
        RECT  17.880 1.360 18.280 1.760 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.780 2.090 ;
        RECT  1.780 1.850 2.310 2.090 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.070 1.690 4.540 2.100 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.710 2.070 0.860 2.470 ;
        RECT  0.860 2.070 1.110 2.650 ;
        RECT  1.110 2.390 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.880 5.440 ;
        RECT  0.880 4.480 1.280 5.440 ;
        RECT  1.280 4.640 4.030 5.440 ;
        RECT  4.030 4.480 4.430 5.440 ;
        RECT  4.430 4.640 6.940 5.440 ;
        RECT  6.940 4.480 7.920 5.440 ;
        RECT  7.920 4.640 14.780 5.440 ;
        RECT  14.780 4.480 15.180 5.440 ;
        RECT  15.180 4.640 16.900 5.440 ;
        RECT  16.900 4.290 16.910 5.440 ;
        RECT  16.910 4.090 17.310 5.440 ;
        RECT  17.310 4.290 17.320 5.440 ;
        RECT  17.320 4.640 19.140 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 2.370 0.400 ;
        RECT  2.370 -0.400 2.770 0.560 ;
        RECT  2.770 -0.400 4.400 0.400 ;
        RECT  4.400 -0.400 4.800 0.560 ;
        RECT  4.800 -0.400 7.360 0.400 ;
        RECT  7.360 -0.400 7.370 1.160 ;
        RECT  7.370 -0.400 7.770 1.360 ;
        RECT  7.770 -0.400 7.780 1.160 ;
        RECT  7.780 -0.400 13.140 0.400 ;
        RECT  13.140 -0.400 13.540 0.560 ;
        RECT  13.540 -0.400 15.910 0.400 ;
        RECT  15.910 -0.400 16.310 0.560 ;
        RECT  16.310 -0.400 17.250 0.400 ;
        RECT  17.250 -0.400 17.260 0.880 ;
        RECT  17.260 -0.400 17.660 1.080 ;
        RECT  17.660 -0.400 17.670 0.880 ;
        RECT  17.670 -0.400 19.140 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  18.130 2.180 18.370 3.780 ;
        RECT  17.890 2.180 18.130 2.580 ;
        RECT  15.980 3.540 18.130 3.780 ;
        RECT  15.950 3.540 15.980 4.180 ;
        RECT  15.720 1.350 15.950 4.180 ;
        RECT  15.710 1.190 15.720 4.180 ;
        RECT  15.320 1.190 15.710 1.590 ;
        RECT  15.580 3.540 15.710 4.180 ;
        RECT  13.640 3.940 15.580 4.180 ;
        RECT  15.260 2.080 15.380 2.480 ;
        RECT  15.020 1.870 15.260 3.660 ;
        RECT  14.980 1.870 15.020 2.110 ;
        RECT  13.960 3.420 15.020 3.660 ;
        RECT  14.740 1.330 14.980 2.110 ;
        RECT  14.580 1.330 14.740 1.730 ;
        RECT  14.340 2.390 14.740 2.790 ;
        RECT  13.360 1.490 14.580 1.730 ;
        RECT  13.120 2.420 14.340 2.790 ;
        RECT  13.400 3.940 13.640 4.360 ;
        RECT  8.430 4.120 13.400 4.360 ;
        RECT  13.120 1.490 13.360 2.140 ;
        RECT  12.880 2.420 13.120 3.760 ;
        RECT  12.840 2.420 12.880 2.660 ;
        RECT  11.960 3.520 12.880 3.760 ;
        RECT  12.600 1.390 12.840 2.660 ;
        RECT  12.340 1.390 12.600 1.630 ;
        RECT  12.320 2.950 12.600 3.190 ;
        RECT  12.100 1.190 12.340 1.630 ;
        RECT  12.080 1.910 12.320 3.190 ;
        RECT  11.680 1.190 12.100 1.430 ;
        RECT  11.820 1.910 12.080 2.150 ;
        RECT  11.430 1.790 11.820 2.150 ;
        RECT  11.680 2.430 11.800 2.830 ;
        RECT  11.440 2.430 11.680 3.830 ;
        RECT  10.670 2.430 11.440 2.670 ;
        RECT  8.950 3.590 11.440 3.830 ;
        RECT  11.190 1.790 11.430 2.030 ;
        RECT  10.950 1.190 11.190 2.030 ;
        RECT  10.750 2.950 11.150 3.310 ;
        RECT  9.860 1.190 10.950 1.430 ;
        RECT  9.470 3.070 10.750 3.310 ;
        RECT  10.430 1.710 10.670 2.670 ;
        RECT  10.340 1.710 10.430 2.110 ;
        RECT  9.990 2.550 10.150 2.790 ;
        RECT  9.860 1.760 9.990 2.790 ;
        RECT  9.750 1.190 9.860 2.790 ;
        RECT  9.620 1.190 9.750 2.080 ;
        RECT  9.340 2.810 9.470 3.310 ;
        RECT  9.230 1.190 9.340 3.310 ;
        RECT  9.100 1.190 9.230 3.050 ;
        RECT  8.800 1.190 9.100 1.430 ;
        RECT  7.740 2.810 9.100 3.050 ;
        RECT  8.710 3.420 8.950 3.830 ;
        RECT  8.580 1.710 8.820 2.410 ;
        RECT  6.940 3.420 8.710 3.660 ;
        RECT  7.460 2.170 8.580 2.410 ;
        RECT  8.190 3.940 8.430 4.360 ;
        RECT  3.590 3.940 8.190 4.180 ;
        RECT  7.420 2.690 7.740 3.050 ;
        RECT  7.220 2.030 7.460 2.410 ;
        RECT  7.340 2.690 7.420 2.930 ;
        RECT  6.370 2.030 7.220 2.270 ;
        RECT  6.700 2.610 6.940 3.660 ;
        RECT  5.770 3.420 6.700 3.660 ;
        RECT  6.370 1.010 6.430 1.410 ;
        RECT  6.130 1.010 6.370 3.140 ;
        RECT  6.030 1.010 6.130 1.410 ;
        RECT  5.750 1.680 5.770 3.660 ;
        RECT  5.530 1.570 5.750 3.660 ;
        RECT  3.510 1.050 5.550 1.290 ;
        RECT  5.350 1.570 5.530 1.970 ;
        RECT  2.890 2.890 5.530 3.130 ;
        RECT  2.830 2.370 5.250 2.610 ;
        RECT  3.170 3.400 5.110 3.640 ;
        RECT  3.170 3.940 3.590 4.220 ;
        RECT  3.110 1.000 3.510 1.400 ;
        RECT  2.610 3.980 3.170 4.220 ;
        RECT  2.650 2.890 2.890 3.670 ;
        RECT  2.590 1.230 2.830 2.610 ;
        RECT  0.490 3.430 2.650 3.670 ;
        RECT  1.710 1.230 2.590 1.470 ;
        RECT  2.370 2.370 2.590 2.610 ;
        RECT  2.130 2.370 2.370 3.150 ;
        RECT  0.410 1.160 0.570 1.560 ;
        RECT  0.410 2.800 0.490 3.670 ;
        RECT  0.250 1.160 0.410 3.670 ;
        RECT  0.170 1.160 0.250 3.190 ;
    END
END JKFFSX2

MACRO JKFFSX1
    CLASS CORE ;
    FOREIGN JKFFSX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFSXL ;
    SIZE 17.820 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.780 1.650 8.050 1.890 ;
        RECT  8.050 0.670 8.290 1.890 ;
        RECT  8.290 0.670 12.620 0.910 ;
        RECT  12.620 0.670 12.860 1.100 ;
        RECT  12.860 0.860 13.820 1.100 ;
        RECT  13.820 0.670 14.220 1.100 ;
        RECT  14.220 0.710 14.320 0.970 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.600 2.970 15.880 3.410 ;
        RECT  15.600 1.390 15.880 1.790 ;
        RECT  15.880 1.390 16.000 3.410 ;
        RECT  16.000 1.470 16.120 3.210 ;
        RECT  16.120 2.950 16.300 3.210 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.250 2.950 17.370 3.350 ;
        RECT  17.360 2.390 17.370 2.650 ;
        RECT  17.250 1.320 17.370 1.960 ;
        RECT  17.370 1.320 17.610 3.350 ;
        RECT  17.610 2.390 17.620 2.650 ;
        RECT  17.610 2.950 17.650 3.350 ;
        RECT  17.610 1.320 17.650 1.960 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.780 2.090 ;
        RECT  1.780 1.850 2.310 2.090 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.070 1.690 4.540 2.100 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.710 2.070 0.860 2.470 ;
        RECT  0.860 2.070 1.110 2.650 ;
        RECT  1.110 2.390 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.880 5.440 ;
        RECT  0.880 4.480 1.280 5.440 ;
        RECT  1.280 4.640 4.030 5.440 ;
        RECT  4.030 4.480 4.430 5.440 ;
        RECT  4.430 4.640 6.940 5.440 ;
        RECT  6.940 4.480 7.920 5.440 ;
        RECT  7.920 4.640 14.200 5.440 ;
        RECT  14.200 4.480 15.180 5.440 ;
        RECT  15.180 4.640 16.420 5.440 ;
        RECT  16.420 4.480 16.820 5.440 ;
        RECT  16.820 4.640 17.820 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 2.370 0.400 ;
        RECT  2.370 -0.400 2.770 0.560 ;
        RECT  2.770 -0.400 4.400 0.400 ;
        RECT  4.400 -0.400 4.800 0.560 ;
        RECT  4.800 -0.400 7.360 0.400 ;
        RECT  7.360 -0.400 7.370 1.160 ;
        RECT  7.370 -0.400 7.770 1.360 ;
        RECT  7.770 -0.400 7.780 1.160 ;
        RECT  7.780 -0.400 13.140 0.400 ;
        RECT  13.140 -0.400 13.540 0.560 ;
        RECT  13.540 -0.400 16.430 0.400 ;
        RECT  16.430 -0.400 16.830 0.560 ;
        RECT  16.830 -0.400 17.820 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.970 2.190 17.000 2.590 ;
        RECT  16.730 0.860 16.970 4.180 ;
        RECT  16.000 0.860 16.730 1.100 ;
        RECT  16.000 3.940 16.730 4.180 ;
        RECT  15.600 0.670 16.000 1.100 ;
        RECT  15.600 3.940 16.000 4.350 ;
        RECT  13.640 3.940 15.600 4.180 ;
        RECT  15.180 2.130 15.380 2.530 ;
        RECT  14.940 1.330 15.180 3.660 ;
        RECT  14.780 1.330 14.940 1.730 ;
        RECT  13.990 3.420 14.940 3.660 ;
        RECT  13.360 1.490 14.780 1.730 ;
        RECT  13.120 2.650 14.660 3.050 ;
        RECT  13.400 3.940 13.640 4.360 ;
        RECT  8.430 4.120 13.400 4.360 ;
        RECT  13.120 1.490 13.360 2.140 ;
        RECT  12.880 2.430 13.120 3.760 ;
        RECT  12.840 2.430 12.880 2.670 ;
        RECT  11.960 3.520 12.880 3.760 ;
        RECT  12.600 1.390 12.840 2.670 ;
        RECT  12.340 1.390 12.600 1.630 ;
        RECT  12.320 2.950 12.600 3.190 ;
        RECT  12.100 1.190 12.340 1.630 ;
        RECT  12.080 1.910 12.320 3.190 ;
        RECT  11.680 1.190 12.100 1.430 ;
        RECT  11.820 1.910 12.080 2.150 ;
        RECT  11.430 1.790 11.820 2.150 ;
        RECT  11.680 2.430 11.800 2.830 ;
        RECT  11.440 2.430 11.680 3.830 ;
        RECT  10.670 2.430 11.440 2.670 ;
        RECT  8.950 3.590 11.440 3.830 ;
        RECT  11.190 1.790 11.430 2.030 ;
        RECT  10.950 1.190 11.190 2.030 ;
        RECT  11.070 2.950 11.150 3.190 ;
        RECT  10.750 2.950 11.070 3.310 ;
        RECT  9.860 1.190 10.950 1.430 ;
        RECT  9.470 3.070 10.750 3.310 ;
        RECT  10.580 1.790 10.670 2.670 ;
        RECT  10.430 1.710 10.580 2.670 ;
        RECT  10.340 1.710 10.430 2.110 ;
        RECT  9.990 2.550 10.150 2.790 ;
        RECT  9.860 1.760 9.990 2.790 ;
        RECT  9.750 1.190 9.860 2.790 ;
        RECT  9.620 1.190 9.750 2.080 ;
        RECT  9.340 2.810 9.470 3.310 ;
        RECT  9.230 1.190 9.340 3.310 ;
        RECT  9.100 1.190 9.230 3.050 ;
        RECT  8.800 1.190 9.100 1.430 ;
        RECT  7.740 2.810 9.100 3.050 ;
        RECT  8.710 3.420 8.950 3.830 ;
        RECT  8.580 1.710 8.820 2.410 ;
        RECT  6.940 3.420 8.710 3.660 ;
        RECT  7.460 2.170 8.580 2.410 ;
        RECT  8.190 3.940 8.430 4.360 ;
        RECT  3.590 3.940 8.190 4.180 ;
        RECT  7.420 2.690 7.740 3.050 ;
        RECT  7.220 2.030 7.460 2.410 ;
        RECT  7.340 2.690 7.420 2.930 ;
        RECT  6.370 2.030 7.220 2.270 ;
        RECT  6.700 2.610 6.940 3.660 ;
        RECT  5.770 3.420 6.700 3.660 ;
        RECT  6.370 1.010 6.430 1.410 ;
        RECT  6.130 1.010 6.370 3.140 ;
        RECT  6.030 1.010 6.130 1.410 ;
        RECT  5.750 1.680 5.770 3.660 ;
        RECT  5.530 1.570 5.750 3.660 ;
        RECT  3.510 1.050 5.550 1.290 ;
        RECT  5.350 1.570 5.530 1.970 ;
        RECT  2.890 2.890 5.530 3.130 ;
        RECT  2.830 2.370 5.250 2.610 ;
        RECT  3.170 3.400 5.110 3.640 ;
        RECT  3.170 3.940 3.590 4.220 ;
        RECT  3.110 1.000 3.510 1.400 ;
        RECT  2.610 3.980 3.170 4.220 ;
        RECT  2.650 2.890 2.890 3.670 ;
        RECT  2.590 1.230 2.830 2.610 ;
        RECT  0.490 3.430 2.650 3.670 ;
        RECT  1.710 1.230 2.590 1.470 ;
        RECT  2.370 2.370 2.590 2.610 ;
        RECT  2.130 2.370 2.370 3.150 ;
        RECT  0.410 1.220 0.570 1.620 ;
        RECT  0.410 2.800 0.490 3.670 ;
        RECT  0.250 1.220 0.410 3.670 ;
        RECT  0.170 1.220 0.250 3.190 ;
    END
END JKFFSX1

MACRO JKFFRXL
    CLASS CORE ;
    FOREIGN JKFFRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.800 1.800 10.450 2.100 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.870 2.980 16.900 3.380 ;
        RECT  16.700 1.270 16.900 1.530 ;
        RECT  16.900 0.860 17.140 3.380 ;
        RECT  17.140 0.860 17.370 1.100 ;
        RECT  17.370 0.710 17.770 1.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.020 2.950 18.130 3.210 ;
        RECT  18.130 2.940 18.430 3.220 ;
        RECT  18.430 2.940 18.570 3.350 ;
        RECT  18.290 1.390 18.570 1.790 ;
        RECT  18.570 1.390 18.690 3.350 ;
        RECT  18.690 1.550 18.810 3.350 ;
        RECT  18.810 2.950 18.830 3.350 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.530 2.090 ;
        RECT  1.530 1.810 1.780 2.090 ;
        RECT  1.780 1.810 2.260 2.050 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 1.270 4.170 1.530 ;
        RECT  4.170 1.270 4.420 1.980 ;
        RECT  4.420 1.530 4.510 1.980 ;
        RECT  4.510 1.580 4.570 1.980 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.720 2.050 0.770 2.450 ;
        RECT  0.770 2.040 1.120 2.660 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.780 5.440 ;
        RECT  0.780 4.480 1.180 5.440 ;
        RECT  1.180 4.640 4.050 5.440 ;
        RECT  4.050 4.480 4.450 5.440 ;
        RECT  4.450 4.640 7.450 5.440 ;
        RECT  7.450 4.480 8.990 5.440 ;
        RECT  8.990 4.640 14.560 5.440 ;
        RECT  14.560 4.480 14.960 5.440 ;
        RECT  14.960 4.640 17.610 5.440 ;
        RECT  17.610 4.480 18.010 5.440 ;
        RECT  18.010 4.640 19.140 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 2.580 0.400 ;
        RECT  2.580 -0.400 2.980 0.560 ;
        RECT  2.980 -0.400 7.460 0.400 ;
        RECT  7.460 -0.400 7.470 1.040 ;
        RECT  7.470 -0.400 7.870 1.240 ;
        RECT  7.870 -0.400 7.880 1.040 ;
        RECT  7.880 -0.400 9.220 0.400 ;
        RECT  9.220 -0.400 9.230 0.810 ;
        RECT  9.230 -0.400 9.630 1.010 ;
        RECT  9.630 -0.400 9.640 0.810 ;
        RECT  9.640 -0.400 14.020 0.400 ;
        RECT  14.020 -0.400 15.000 0.560 ;
        RECT  15.000 -0.400 16.490 0.400 ;
        RECT  16.490 -0.400 16.890 0.560 ;
        RECT  16.890 -0.400 18.260 0.400 ;
        RECT  18.260 -0.400 18.660 0.560 ;
        RECT  18.660 -0.400 19.140 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  17.690 2.130 18.330 2.530 ;
        RECT  17.660 1.390 17.690 2.530 ;
        RECT  17.450 1.390 17.660 4.040 ;
        RECT  17.420 2.290 17.450 4.040 ;
        RECT  17.050 3.800 17.420 4.040 ;
        RECT  16.810 3.800 17.050 4.280 ;
        RECT  15.470 4.040 16.810 4.280 ;
        RECT  16.500 2.300 16.620 2.700 ;
        RECT  16.260 1.810 16.500 3.760 ;
        RECT  16.120 1.810 16.260 2.050 ;
        RECT  15.840 3.520 16.260 3.760 ;
        RECT  15.830 1.370 16.120 2.050 ;
        RECT  15.580 2.810 15.980 3.210 ;
        RECT  15.720 1.370 15.830 2.040 ;
        RECT  15.420 0.690 15.820 1.100 ;
        RECT  14.650 1.640 15.720 2.040 ;
        RECT  14.480 2.890 15.580 3.130 ;
        RECT  15.230 3.940 15.470 4.280 ;
        RECT  12.160 0.860 15.420 1.100 ;
        RECT  13.430 3.940 15.230 4.180 ;
        RECT  14.370 2.320 14.480 3.660 ;
        RECT  14.240 1.380 14.370 3.660 ;
        RECT  14.130 1.380 14.240 2.560 ;
        RECT  13.190 3.420 14.240 3.660 ;
        RECT  13.630 1.380 14.130 1.780 ;
        RECT  13.800 2.850 13.960 3.090 ;
        RECT  13.560 2.200 13.800 3.090 ;
        RECT  13.300 2.200 13.560 2.440 ;
        RECT  13.190 3.940 13.430 4.360 ;
        RECT  13.060 1.420 13.300 2.440 ;
        RECT  12.910 2.750 13.240 2.990 ;
        RECT  9.510 4.120 13.190 4.360 ;
        RECT  11.640 1.420 13.060 1.660 ;
        RECT  12.660 2.750 12.910 3.840 ;
        RECT  10.040 3.600 12.660 3.840 ;
        RECT  12.220 2.670 12.380 3.070 ;
        RECT  11.980 2.670 12.220 3.320 ;
        RECT  11.920 0.680 12.160 1.100 ;
        RECT  10.560 3.080 11.980 3.320 ;
        RECT  10.730 0.680 11.920 0.920 ;
        RECT  11.240 1.200 11.640 1.660 ;
        RECT  11.080 1.420 11.240 1.660 ;
        RECT  11.080 2.560 11.240 2.800 ;
        RECT  10.840 1.420 11.080 2.800 ;
        RECT  10.720 1.420 10.840 1.820 ;
        RECT  10.490 0.680 10.730 1.130 ;
        RECT  10.320 2.900 10.560 3.320 ;
        RECT  10.310 0.890 10.490 1.130 ;
        RECT  8.600 2.900 10.320 3.140 ;
        RECT  10.070 0.890 10.310 1.530 ;
        RECT  9.270 2.380 10.280 2.620 ;
        RECT  9.280 1.290 10.070 1.530 ;
        RECT  9.800 3.420 10.040 3.840 ;
        RECT  5.850 3.420 9.800 3.660 ;
        RECT  9.270 3.940 9.510 4.360 ;
        RECT  9.270 1.290 9.280 2.090 ;
        RECT  9.040 1.290 9.270 2.620 ;
        RECT  3.730 3.940 9.270 4.180 ;
        RECT  9.030 1.690 9.040 2.620 ;
        RECT  8.880 1.690 9.030 2.090 ;
        RECT  8.590 0.950 8.750 1.350 ;
        RECT  8.590 2.540 8.600 3.140 ;
        RECT  8.350 0.950 8.590 3.140 ;
        RECT  7.980 2.400 8.350 3.140 ;
        RECT  7.640 1.520 8.040 1.920 ;
        RECT  7.550 2.400 7.980 2.640 ;
        RECT  6.530 1.600 7.640 1.840 ;
        RECT  7.150 2.240 7.550 2.640 ;
        RECT  6.380 1.070 6.530 1.840 ;
        RECT  6.140 1.070 6.380 3.140 ;
        RECT  6.130 1.070 6.140 1.470 ;
        RECT  5.610 1.530 5.850 3.660 ;
        RECT  5.490 1.010 5.650 1.250 ;
        RECT  5.450 1.530 5.610 1.930 ;
        RECT  2.900 2.850 5.610 3.090 ;
        RECT  5.250 0.750 5.490 1.250 ;
        RECT  2.780 2.330 5.330 2.570 ;
        RECT  3.570 0.750 5.250 0.990 ;
        RECT  3.180 3.370 5.120 3.610 ;
        RECT  3.410 3.940 3.730 4.200 ;
        RECT  3.330 0.750 3.570 1.410 ;
        RECT  1.460 3.960 3.410 4.200 ;
        RECT  3.170 1.010 3.330 1.410 ;
        RECT  2.660 2.850 2.900 3.680 ;
        RECT  2.540 1.290 2.780 2.570 ;
        RECT  0.490 3.440 2.660 3.680 ;
        RECT  2.110 1.290 2.540 1.530 ;
        RECT  2.380 2.330 2.540 2.570 ;
        RECT  2.140 2.330 2.380 3.150 ;
        RECT  1.710 1.130 2.110 1.530 ;
        RECT  0.400 1.130 0.570 1.530 ;
        RECT  0.400 2.800 0.490 3.680 ;
        RECT  0.250 1.130 0.400 3.680 ;
        RECT  0.160 1.130 0.250 3.200 ;
    END
END JKFFRXL

MACRO JKFFRX4
    CLASS CORE ;
    FOREIGN JKFFRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFRXL ;
    SIZE 23.760 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.550 1.860 10.100 2.100 ;
        RECT  10.100 1.830 10.360 2.100 ;
        RECT  10.360 1.860 10.530 2.100 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.080 2.830 21.230 3.230 ;
        RECT  21.200 1.150 21.230 1.550 ;
        RECT  21.230 1.150 21.630 3.230 ;
        RECT  21.630 1.150 21.640 2.660 ;
        RECT  21.640 1.260 21.670 2.660 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  22.540 2.830 22.550 3.230 ;
        RECT  22.490 1.150 22.550 1.550 ;
        RECT  22.550 1.150 22.950 3.230 ;
        RECT  22.950 1.260 22.990 2.660 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.530 2.090 ;
        RECT  1.530 1.810 1.780 2.090 ;
        RECT  1.780 1.810 2.420 2.050 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 1.270 4.170 1.530 ;
        RECT  4.170 1.270 4.190 1.850 ;
        RECT  4.190 1.270 4.420 1.930 ;
        RECT  4.420 1.530 4.590 1.930 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.720 2.050 0.770 2.450 ;
        RECT  0.770 2.040 1.120 2.660 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.780 5.440 ;
        RECT  0.780 4.480 1.180 5.440 ;
        RECT  1.180 4.640 4.050 5.440 ;
        RECT  4.050 4.480 4.450 5.440 ;
        RECT  4.450 4.640 7.170 5.440 ;
        RECT  7.170 4.480 8.150 5.440 ;
        RECT  8.150 4.640 14.440 5.440 ;
        RECT  14.440 4.480 14.840 5.440 ;
        RECT  14.840 4.640 16.330 5.440 ;
        RECT  16.330 4.480 16.730 5.440 ;
        RECT  16.730 4.640 18.970 5.440 ;
        RECT  18.970 4.480 19.370 5.440 ;
        RECT  19.370 4.640 20.400 5.440 ;
        RECT  20.400 4.230 20.410 5.440 ;
        RECT  20.410 4.030 20.810 5.440 ;
        RECT  20.810 4.230 20.820 5.440 ;
        RECT  20.820 4.640 21.790 5.440 ;
        RECT  21.790 4.230 21.800 5.440 ;
        RECT  21.800 4.030 22.200 5.440 ;
        RECT  22.200 4.230 22.210 5.440 ;
        RECT  22.210 4.640 23.180 5.440 ;
        RECT  23.180 4.230 23.190 5.440 ;
        RECT  23.190 4.030 23.590 5.440 ;
        RECT  23.590 4.230 23.600 5.440 ;
        RECT  23.600 4.640 23.760 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.830 0.400 ;
        RECT  0.830 -0.400 1.230 0.560 ;
        RECT  1.230 -0.400 2.590 0.400 ;
        RECT  2.590 -0.400 2.990 0.560 ;
        RECT  2.990 -0.400 7.460 0.400 ;
        RECT  7.460 -0.400 7.470 1.110 ;
        RECT  7.470 -0.400 7.870 1.310 ;
        RECT  7.870 -0.400 7.880 1.110 ;
        RECT  7.880 -0.400 9.040 0.400 ;
        RECT  9.040 -0.400 9.050 0.810 ;
        RECT  9.050 -0.400 9.450 1.010 ;
        RECT  9.450 -0.400 9.460 0.810 ;
        RECT  9.460 -0.400 12.510 0.400 ;
        RECT  12.510 -0.400 12.750 1.310 ;
        RECT  12.750 -0.400 14.990 0.400 ;
        RECT  14.990 -0.400 15.390 0.560 ;
        RECT  15.390 -0.400 16.990 0.400 ;
        RECT  16.990 -0.400 17.000 0.730 ;
        RECT  17.000 -0.400 17.400 0.930 ;
        RECT  17.400 -0.400 17.410 0.730 ;
        RECT  17.410 -0.400 18.510 0.400 ;
        RECT  18.510 -0.400 18.520 1.060 ;
        RECT  18.520 -0.400 18.920 1.260 ;
        RECT  18.920 -0.400 18.930 1.060 ;
        RECT  18.930 -0.400 20.510 0.400 ;
        RECT  20.510 -0.400 20.520 0.670 ;
        RECT  20.520 -0.400 20.920 0.870 ;
        RECT  20.920 -0.400 20.930 0.670 ;
        RECT  20.930 -0.400 21.810 0.400 ;
        RECT  21.810 -0.400 21.820 0.670 ;
        RECT  21.820 -0.400 22.220 0.870 ;
        RECT  22.220 -0.400 22.230 0.670 ;
        RECT  22.230 -0.400 23.100 0.400 ;
        RECT  23.100 -0.400 23.110 0.670 ;
        RECT  23.110 -0.400 23.510 0.870 ;
        RECT  23.510 -0.400 23.520 0.670 ;
        RECT  23.520 -0.400 23.760 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  23.230 2.260 23.470 3.750 ;
        RECT  20.840 3.510 23.230 3.750 ;
        RECT  20.600 1.420 20.840 3.750 ;
        RECT  20.010 1.420 20.600 1.660 ;
        RECT  20.010 3.230 20.600 3.750 ;
        RECT  19.530 1.940 20.360 2.340 ;
        RECT  19.770 1.020 20.010 1.660 ;
        RECT  19.770 3.230 20.010 4.180 ;
        RECT  19.680 1.020 19.770 1.260 ;
        RECT  14.080 3.940 19.770 4.180 ;
        RECT  19.280 0.860 19.680 1.260 ;
        RECT  19.290 1.540 19.530 3.500 ;
        RECT  18.160 1.540 19.290 1.780 ;
        RECT  18.110 3.260 19.290 3.500 ;
        RECT  18.770 2.060 19.010 2.780 ;
        RECT  17.650 2.060 18.770 2.300 ;
        RECT  17.940 2.580 18.340 2.980 ;
        RECT  17.920 1.050 18.160 1.780 ;
        RECT  17.710 3.260 18.110 3.660 ;
        RECT  17.000 2.740 17.940 2.980 ;
        RECT  17.760 1.050 17.920 1.460 ;
        RECT  16.720 1.220 17.760 1.460 ;
        RECT  17.410 2.060 17.650 2.460 ;
        RECT  17.250 2.220 17.410 2.460 ;
        RECT  16.760 1.740 17.000 3.660 ;
        RECT  16.140 1.740 16.760 1.980 ;
        RECT  13.560 3.420 16.760 3.660 ;
        RECT  16.480 0.690 16.720 1.460 ;
        RECT  15.900 1.380 16.140 1.980 ;
        RECT  16.060 0.670 16.070 0.910 ;
        RECT  15.670 0.670 16.060 1.100 ;
        RECT  15.570 2.470 15.970 2.870 ;
        RECT  13.710 1.380 15.900 1.620 ;
        RECT  13.270 0.860 15.670 1.100 ;
        RECT  15.500 2.470 15.570 2.710 ;
        RECT  15.260 2.110 15.500 2.710 ;
        RECT  11.710 2.110 15.260 2.350 ;
        RECT  14.580 2.830 14.980 3.140 ;
        RECT  12.880 2.900 14.580 3.140 ;
        RECT  13.840 3.940 14.080 4.370 ;
        RECT  8.660 4.130 13.840 4.370 ;
        RECT  13.160 3.420 13.560 3.820 ;
        RECT  13.030 0.860 13.270 1.830 ;
        RECT  12.230 1.590 13.030 1.830 ;
        RECT  12.640 2.900 12.880 3.840 ;
        RECT  9.180 3.600 12.640 3.840 ;
        RECT  12.120 2.750 12.360 3.320 ;
        RECT  11.990 0.680 12.230 1.830 ;
        RECT  9.700 3.080 12.120 3.320 ;
        RECT  10.290 0.680 11.990 0.920 ;
        RECT  11.540 1.210 11.710 2.350 ;
        RECT  11.310 1.210 11.540 2.360 ;
        RECT  11.200 1.690 11.310 2.360 ;
        RECT  10.800 1.690 11.200 2.800 ;
        RECT  9.980 2.380 10.380 2.800 ;
        RECT  10.050 0.680 10.290 1.530 ;
        RECT  9.870 1.120 10.050 1.530 ;
        RECT  9.210 2.380 9.980 2.620 ;
        RECT  9.210 1.290 9.870 1.530 ;
        RECT  9.460 2.900 9.700 3.320 ;
        RECT  8.540 2.900 9.460 3.140 ;
        RECT  8.970 1.290 9.210 2.620 ;
        RECT  8.940 3.420 9.180 3.840 ;
        RECT  8.810 1.690 8.970 2.090 ;
        RECT  5.780 3.420 8.940 3.660 ;
        RECT  8.420 3.940 8.660 4.370 ;
        RECT  8.530 0.920 8.630 1.320 ;
        RECT  8.530 2.540 8.540 3.140 ;
        RECT  8.290 0.920 8.530 3.140 ;
        RECT  3.730 3.940 8.420 4.180 ;
        RECT  8.230 0.920 8.290 1.320 ;
        RECT  7.980 2.400 8.290 3.140 ;
        RECT  6.530 1.600 8.010 1.840 ;
        RECT  7.550 2.400 7.980 2.640 ;
        RECT  7.150 2.240 7.550 2.640 ;
        RECT  6.380 1.060 6.530 1.840 ;
        RECT  6.140 1.060 6.380 3.140 ;
        RECT  6.130 1.060 6.140 1.460 ;
        RECT  5.780 1.530 5.850 1.930 ;
        RECT  5.540 1.530 5.780 3.660 ;
        RECT  5.490 1.010 5.650 1.250 ;
        RECT  5.450 1.530 5.540 1.930 ;
        RECT  2.900 2.850 5.540 3.090 ;
        RECT  5.250 0.750 5.490 1.250 ;
        RECT  2.930 2.330 5.260 2.570 ;
        RECT  3.570 0.750 5.250 0.990 ;
        RECT  3.180 3.370 5.180 3.610 ;
        RECT  3.410 3.940 3.730 4.200 ;
        RECT  3.330 0.750 3.570 1.410 ;
        RECT  1.460 3.960 3.410 4.200 ;
        RECT  3.170 1.010 3.330 1.410 ;
        RECT  2.690 1.300 2.930 2.570 ;
        RECT  2.660 2.850 2.900 3.680 ;
        RECT  2.110 1.300 2.690 1.540 ;
        RECT  2.380 2.330 2.690 2.570 ;
        RECT  0.570 3.440 2.660 3.680 ;
        RECT  2.140 2.330 2.380 3.150 ;
        RECT  1.710 1.140 2.110 1.540 ;
        RECT  0.400 1.130 0.570 1.530 ;
        RECT  0.400 2.930 0.570 3.680 ;
        RECT  0.330 1.130 0.400 3.680 ;
        RECT  0.160 1.130 0.330 3.330 ;
    END
END JKFFRX4

MACRO JKFFRX2
    CLASS CORE ;
    FOREIGN JKFFRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFRXL ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.800 1.800 10.450 2.100 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.840 1.150 17.930 1.550 ;
        RECT  17.920 2.830 18.030 3.230 ;
        RECT  17.930 1.150 18.030 2.100 ;
        RECT  18.030 1.150 18.270 3.230 ;
        RECT  18.270 1.830 18.280 2.090 ;
        RECT  18.270 2.830 18.320 3.230 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.680 1.270 18.810 1.530 ;
        RECT  18.810 1.260 19.080 1.540 ;
        RECT  19.160 2.890 19.400 3.290 ;
        RECT  19.080 1.150 19.400 1.550 ;
        RECT  19.400 1.150 19.480 3.290 ;
        RECT  19.480 1.230 19.560 3.290 ;
        RECT  19.560 1.230 19.640 3.210 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.540 2.090 ;
        RECT  1.540 1.820 1.780 2.090 ;
        RECT  1.780 1.820 1.900 2.060 ;
        RECT  1.900 1.810 2.140 2.060 ;
        RECT  2.140 1.810 2.300 2.050 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 1.270 4.170 1.530 ;
        RECT  4.170 1.270 4.190 1.850 ;
        RECT  4.190 1.270 4.420 1.930 ;
        RECT  4.420 1.530 4.590 1.930 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.720 2.050 0.770 2.450 ;
        RECT  0.770 2.040 1.120 2.660 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.780 5.440 ;
        RECT  0.780 4.480 1.180 5.440 ;
        RECT  1.180 4.640 4.050 5.440 ;
        RECT  4.050 4.480 4.450 5.440 ;
        RECT  4.450 4.640 7.200 5.440 ;
        RECT  7.200 4.480 8.180 5.440 ;
        RECT  8.180 4.640 14.560 5.440 ;
        RECT  14.560 4.480 14.960 5.440 ;
        RECT  14.960 4.640 16.570 5.440 ;
        RECT  16.570 4.480 16.970 5.440 ;
        RECT  16.970 4.640 18.530 5.440 ;
        RECT  18.530 4.230 18.540 5.440 ;
        RECT  18.540 4.030 18.940 5.440 ;
        RECT  18.940 4.230 18.950 5.440 ;
        RECT  18.950 4.640 19.800 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 2.580 0.400 ;
        RECT  2.580 -0.400 2.980 0.560 ;
        RECT  2.980 -0.400 7.460 0.400 ;
        RECT  7.460 -0.400 7.470 1.040 ;
        RECT  7.470 -0.400 7.870 1.240 ;
        RECT  7.870 -0.400 7.880 1.040 ;
        RECT  7.880 -0.400 9.220 0.400 ;
        RECT  9.220 -0.400 9.230 0.810 ;
        RECT  9.230 -0.400 9.630 1.010 ;
        RECT  9.630 -0.400 9.640 0.810 ;
        RECT  9.640 -0.400 13.510 0.400 ;
        RECT  13.510 -0.400 15.050 0.560 ;
        RECT  15.050 -0.400 16.330 0.400 ;
        RECT  16.330 -0.400 16.340 1.360 ;
        RECT  16.340 -0.400 16.740 1.560 ;
        RECT  16.740 -0.400 16.750 1.360 ;
        RECT  16.750 -0.400 18.450 0.400 ;
        RECT  18.450 -0.400 18.460 0.670 ;
        RECT  18.460 -0.400 18.860 0.870 ;
        RECT  18.860 -0.400 18.870 0.670 ;
        RECT  18.870 -0.400 19.800 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  18.880 1.830 19.120 2.610 ;
        RECT  18.840 2.370 18.880 2.610 ;
        RECT  18.600 2.370 18.840 3.750 ;
        RECT  17.580 3.510 18.600 3.750 ;
        RECT  17.420 3.080 17.580 3.750 ;
        RECT  17.420 1.300 17.500 1.700 ;
        RECT  17.180 1.300 17.420 4.180 ;
        RECT  17.100 1.300 17.180 1.700 ;
        RECT  14.270 3.940 17.180 4.180 ;
        RECT  16.700 2.070 16.860 3.470 ;
        RECT  16.460 1.940 16.700 3.470 ;
        RECT  15.990 1.940 16.460 2.180 ;
        RECT  16.240 3.150 16.460 3.470 ;
        RECT  15.840 3.150 16.240 3.550 ;
        RECT  15.780 2.460 16.180 2.860 ;
        RECT  15.980 1.500 15.990 2.180 ;
        RECT  15.650 1.380 15.980 2.180 ;
        RECT  14.480 2.540 15.780 2.780 ;
        RECT  15.340 0.670 15.740 1.100 ;
        RECT  15.580 1.380 15.650 2.000 ;
        RECT  15.570 1.500 15.580 2.000 ;
        RECT  14.690 1.580 15.570 2.000 ;
        RECT  11.810 0.860 15.340 1.100 ;
        RECT  14.570 1.590 14.690 1.990 ;
        RECT  14.280 2.320 14.480 3.660 ;
        RECT  14.240 1.380 14.280 3.660 ;
        RECT  14.030 3.940 14.270 4.360 ;
        RECT  14.040 1.380 14.240 2.560 ;
        RECT  13.590 3.420 14.240 3.660 ;
        RECT  13.300 1.380 14.040 1.780 ;
        RECT  8.690 4.120 14.030 4.360 ;
        RECT  13.760 2.900 13.960 3.140 ;
        RECT  13.520 2.200 13.760 3.140 ;
        RECT  13.190 3.420 13.590 3.840 ;
        RECT  12.970 2.200 13.520 2.440 ;
        RECT  12.910 2.830 13.240 3.070 ;
        RECT  12.730 1.420 12.970 2.440 ;
        RECT  12.660 2.830 12.910 3.840 ;
        RECT  11.290 1.420 12.730 1.660 ;
        RECT  9.210 3.600 12.660 3.840 ;
        RECT  11.980 2.750 12.380 3.320 ;
        RECT  9.730 3.080 11.980 3.320 ;
        RECT  11.570 0.680 11.810 1.100 ;
        RECT  10.450 0.680 11.570 0.920 ;
        RECT  11.040 1.200 11.290 1.660 ;
        RECT  11.040 2.560 11.200 2.800 ;
        RECT  10.800 1.200 11.040 2.800 ;
        RECT  10.720 1.690 10.800 2.090 ;
        RECT  10.060 2.380 10.460 2.800 ;
        RECT  10.290 0.680 10.450 1.320 ;
        RECT  10.050 0.680 10.290 1.530 ;
        RECT  9.270 2.380 10.060 2.620 ;
        RECT  9.280 1.290 10.050 1.530 ;
        RECT  9.490 2.900 9.730 3.320 ;
        RECT  8.600 2.900 9.490 3.140 ;
        RECT  9.270 1.290 9.280 2.090 ;
        RECT  9.040 1.290 9.270 2.620 ;
        RECT  8.970 3.420 9.210 3.840 ;
        RECT  9.030 1.690 9.040 2.620 ;
        RECT  8.880 1.690 9.030 2.090 ;
        RECT  5.780 3.420 8.970 3.660 ;
        RECT  8.590 0.960 8.750 1.360 ;
        RECT  8.450 3.940 8.690 4.360 ;
        RECT  8.590 2.540 8.600 3.140 ;
        RECT  8.350 0.960 8.590 3.140 ;
        RECT  3.730 3.940 8.450 4.180 ;
        RECT  7.980 2.400 8.350 3.140 ;
        RECT  7.640 1.520 8.040 1.920 ;
        RECT  7.550 2.400 7.980 2.640 ;
        RECT  6.530 1.600 7.640 1.840 ;
        RECT  7.150 2.240 7.550 2.640 ;
        RECT  6.380 1.070 6.530 1.840 ;
        RECT  6.140 1.070 6.380 3.140 ;
        RECT  6.130 1.070 6.140 1.470 ;
        RECT  5.780 1.530 5.850 1.930 ;
        RECT  5.540 1.530 5.780 3.660 ;
        RECT  5.490 1.010 5.650 1.250 ;
        RECT  5.450 1.530 5.540 1.930 ;
        RECT  2.900 2.850 5.540 3.090 ;
        RECT  5.250 0.750 5.490 1.250 ;
        RECT  2.780 2.330 5.260 2.570 ;
        RECT  3.570 0.750 5.250 0.990 ;
        RECT  3.180 3.360 5.120 3.600 ;
        RECT  3.410 3.940 3.730 4.200 ;
        RECT  3.330 0.750 3.570 1.410 ;
        RECT  1.460 3.960 3.410 4.200 ;
        RECT  3.170 1.010 3.330 1.410 ;
        RECT  2.660 2.850 2.900 3.680 ;
        RECT  2.540 1.300 2.780 2.570 ;
        RECT  0.490 3.440 2.660 3.680 ;
        RECT  2.110 1.300 2.540 1.540 ;
        RECT  2.380 2.330 2.540 2.570 ;
        RECT  2.140 2.330 2.380 3.150 ;
        RECT  1.710 1.140 2.110 1.540 ;
        RECT  0.400 1.130 0.570 1.530 ;
        RECT  0.400 2.800 0.490 3.680 ;
        RECT  0.250 1.130 0.400 3.680 ;
        RECT  0.160 1.130 0.250 3.200 ;
    END
END JKFFRX2

MACRO JKFFRX1
    CLASS CORE ;
    FOREIGN JKFFRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFRXL ;
    SIZE 19.140 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.800 1.800 10.450 2.100 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.870 2.980 16.900 3.380 ;
        RECT  16.700 1.270 16.900 1.530 ;
        RECT  16.900 0.860 17.140 3.380 ;
        RECT  17.140 0.860 17.310 1.100 ;
        RECT  17.310 0.710 17.720 1.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.020 2.950 18.130 3.210 ;
        RECT  18.130 2.940 18.430 3.220 ;
        RECT  18.430 2.940 18.570 3.350 ;
        RECT  18.350 1.320 18.570 1.720 ;
        RECT  18.570 1.320 18.750 3.350 ;
        RECT  18.750 1.480 18.810 3.350 ;
        RECT  18.810 2.950 18.830 3.350 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.540 2.090 ;
        RECT  1.540 1.820 1.780 2.090 ;
        RECT  1.780 1.820 1.900 2.060 ;
        RECT  1.900 1.770 2.140 2.060 ;
        RECT  2.140 1.770 2.300 2.010 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 1.270 4.170 1.530 ;
        RECT  4.170 1.270 4.190 1.850 ;
        RECT  4.190 1.270 4.420 1.930 ;
        RECT  4.420 1.530 4.590 1.930 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.720 2.050 0.770 2.450 ;
        RECT  0.770 2.040 1.120 2.660 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.780 5.440 ;
        RECT  0.780 4.480 1.180 5.440 ;
        RECT  1.180 4.640 4.050 5.440 ;
        RECT  4.050 4.480 4.450 5.440 ;
        RECT  4.450 4.640 7.450 5.440 ;
        RECT  7.450 4.480 8.990 5.440 ;
        RECT  8.990 4.640 14.560 5.440 ;
        RECT  14.560 4.480 14.960 5.440 ;
        RECT  14.960 4.640 17.610 5.440 ;
        RECT  17.610 4.480 18.010 5.440 ;
        RECT  18.010 4.640 19.140 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 2.580 0.400 ;
        RECT  2.580 -0.400 2.980 0.560 ;
        RECT  2.980 -0.400 7.460 0.400 ;
        RECT  7.460 -0.400 7.470 1.040 ;
        RECT  7.470 -0.400 7.870 1.240 ;
        RECT  7.870 -0.400 7.880 1.040 ;
        RECT  7.880 -0.400 9.220 0.400 ;
        RECT  9.220 -0.400 9.230 0.810 ;
        RECT  9.230 -0.400 9.630 1.010 ;
        RECT  9.630 -0.400 9.640 0.810 ;
        RECT  9.640 -0.400 13.660 0.400 ;
        RECT  13.660 -0.400 15.200 0.560 ;
        RECT  15.200 -0.400 16.490 0.400 ;
        RECT  16.490 -0.400 16.890 0.560 ;
        RECT  16.890 -0.400 18.210 0.400 ;
        RECT  18.210 -0.400 18.610 0.560 ;
        RECT  18.610 -0.400 19.140 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  17.690 2.000 18.330 2.400 ;
        RECT  17.660 1.390 17.690 2.400 ;
        RECT  17.450 1.390 17.660 4.180 ;
        RECT  17.420 2.160 17.450 4.180 ;
        RECT  17.190 3.940 17.420 4.180 ;
        RECT  16.790 3.940 17.190 4.340 ;
        RECT  15.470 4.040 16.790 4.280 ;
        RECT  16.500 2.300 16.620 2.700 ;
        RECT  16.260 1.810 16.500 3.760 ;
        RECT  16.070 1.810 16.260 2.050 ;
        RECT  15.840 3.520 16.260 3.760 ;
        RECT  15.830 1.380 16.070 2.050 ;
        RECT  15.580 2.810 15.980 3.210 ;
        RECT  15.470 0.690 15.870 1.100 ;
        RECT  15.670 1.380 15.830 2.040 ;
        RECT  14.650 1.640 15.670 2.040 ;
        RECT  14.480 2.890 15.580 3.130 ;
        RECT  12.160 0.860 15.470 1.100 ;
        RECT  15.230 3.940 15.470 4.280 ;
        RECT  13.430 3.940 15.230 4.180 ;
        RECT  14.370 2.320 14.480 3.660 ;
        RECT  14.240 1.380 14.370 3.660 ;
        RECT  14.130 1.380 14.240 2.560 ;
        RECT  13.190 3.420 14.240 3.660 ;
        RECT  13.630 1.380 14.130 1.780 ;
        RECT  13.800 2.850 13.960 3.090 ;
        RECT  13.560 2.200 13.800 3.090 ;
        RECT  13.300 2.200 13.560 2.440 ;
        RECT  13.190 3.940 13.430 4.360 ;
        RECT  13.060 1.420 13.300 2.440 ;
        RECT  12.910 2.830 13.240 3.070 ;
        RECT  9.510 4.120 13.190 4.360 ;
        RECT  11.640 1.420 13.060 1.660 ;
        RECT  12.660 2.830 12.910 3.840 ;
        RECT  10.040 3.600 12.660 3.840 ;
        RECT  11.980 2.770 12.380 3.320 ;
        RECT  11.920 0.680 12.160 1.100 ;
        RECT  10.560 3.080 11.980 3.320 ;
        RECT  10.730 0.680 11.920 0.920 ;
        RECT  11.240 1.200 11.640 1.660 ;
        RECT  11.080 1.420 11.240 1.660 ;
        RECT  11.080 2.560 11.240 2.800 ;
        RECT  10.840 1.420 11.080 2.800 ;
        RECT  10.720 1.420 10.840 1.820 ;
        RECT  10.490 0.680 10.730 1.130 ;
        RECT  10.320 2.900 10.560 3.320 ;
        RECT  10.310 0.890 10.490 1.130 ;
        RECT  8.600 2.900 10.320 3.140 ;
        RECT  10.070 0.890 10.310 1.530 ;
        RECT  9.270 2.380 10.280 2.620 ;
        RECT  9.280 1.290 10.070 1.530 ;
        RECT  9.800 3.420 10.040 3.840 ;
        RECT  5.780 3.420 9.800 3.660 ;
        RECT  9.270 3.940 9.510 4.360 ;
        RECT  9.270 1.290 9.280 2.090 ;
        RECT  9.040 1.290 9.270 2.620 ;
        RECT  3.730 3.940 9.270 4.180 ;
        RECT  9.030 1.690 9.040 2.620 ;
        RECT  8.880 1.690 9.030 2.090 ;
        RECT  8.590 0.950 8.750 1.350 ;
        RECT  8.590 2.540 8.600 3.140 ;
        RECT  8.350 0.950 8.590 3.140 ;
        RECT  7.980 2.400 8.350 3.140 ;
        RECT  7.640 1.520 8.040 1.920 ;
        RECT  7.550 2.400 7.980 2.640 ;
        RECT  6.530 1.600 7.640 1.840 ;
        RECT  7.150 2.240 7.550 2.640 ;
        RECT  6.380 1.070 6.530 1.840 ;
        RECT  6.140 1.070 6.380 3.140 ;
        RECT  6.130 1.070 6.140 1.470 ;
        RECT  5.780 1.530 5.850 1.930 ;
        RECT  5.540 1.530 5.780 3.660 ;
        RECT  5.490 1.010 5.650 1.250 ;
        RECT  5.450 1.530 5.540 1.930 ;
        RECT  2.900 2.850 5.540 3.090 ;
        RECT  5.250 0.750 5.490 1.250 ;
        RECT  2.780 2.330 5.260 2.570 ;
        RECT  3.570 0.750 5.250 0.990 ;
        RECT  3.180 3.360 5.120 3.600 ;
        RECT  3.410 3.940 3.730 4.200 ;
        RECT  3.330 0.750 3.570 1.410 ;
        RECT  1.460 3.960 3.410 4.200 ;
        RECT  3.170 1.010 3.330 1.410 ;
        RECT  2.660 2.850 2.900 3.680 ;
        RECT  2.540 1.290 2.780 2.570 ;
        RECT  0.490 3.440 2.660 3.680 ;
        RECT  2.110 1.290 2.540 1.530 ;
        RECT  2.380 2.330 2.540 2.570 ;
        RECT  2.140 2.330 2.380 3.150 ;
        RECT  1.710 1.130 2.110 1.530 ;
        RECT  0.400 1.130 0.570 1.530 ;
        RECT  0.400 2.800 0.490 3.680 ;
        RECT  0.250 1.130 0.400 3.680 ;
        RECT  0.160 1.130 0.250 3.200 ;
    END
END JKFFRX1

MACRO JKFFXL
    CLASS CORE ;
    FOREIGN JKFFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.740 2.950 12.940 3.210 ;
        RECT  12.940 2.810 12.990 3.210 ;
        RECT  12.990 1.380 13.230 3.210 ;
        RECT  13.230 2.810 13.340 3.210 ;
        RECT  13.230 1.380 13.390 1.780 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.610 2.840 14.630 3.240 ;
        RECT  14.630 2.570 14.720 3.240 ;
        RECT  14.720 2.390 14.730 3.240 ;
        RECT  14.610 1.400 14.730 1.910 ;
        RECT  14.730 1.400 14.970 3.240 ;
        RECT  14.970 2.390 14.980 3.240 ;
        RECT  14.980 2.570 15.010 3.240 ;
        RECT  14.970 1.400 15.010 1.910 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.510 2.090 ;
        RECT  3.510 1.830 3.760 2.220 ;
        RECT  3.760 1.980 4.160 2.220 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.570 3.500 0.850 3.900 ;
        RECT  0.850 3.490 1.120 3.910 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.810 2.050 2.230 ;
        RECT  2.050 1.820 2.280 2.220 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.750 5.440 ;
        RECT  1.750 3.890 1.760 5.440 ;
        RECT  1.760 3.690 2.160 5.440 ;
        RECT  2.160 3.890 2.170 5.440 ;
        RECT  2.170 4.640 4.190 5.440 ;
        RECT  4.190 4.180 4.200 5.440 ;
        RECT  4.200 4.060 4.600 5.440 ;
        RECT  4.600 4.180 4.610 5.440 ;
        RECT  4.610 4.640 7.190 5.440 ;
        RECT  7.190 3.980 7.430 5.440 ;
        RECT  7.430 4.640 9.180 5.440 ;
        RECT  9.180 3.680 9.190 5.440 ;
        RECT  9.190 3.480 9.590 5.440 ;
        RECT  9.590 3.680 9.600 5.440 ;
        RECT  9.600 4.640 12.120 5.440 ;
        RECT  12.120 4.480 12.520 5.440 ;
        RECT  12.520 4.640 13.780 5.440 ;
        RECT  13.780 4.480 14.180 5.440 ;
        RECT  14.180 4.640 15.180 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.500 0.400 ;
        RECT  1.500 -0.400 1.900 0.560 ;
        RECT  1.900 -0.400 6.390 0.400 ;
        RECT  6.390 -0.400 7.370 0.560 ;
        RECT  7.370 -0.400 8.640 0.400 ;
        RECT  8.640 -0.400 8.650 1.040 ;
        RECT  8.650 -0.400 9.050 1.240 ;
        RECT  9.050 -0.400 9.060 1.040 ;
        RECT  9.060 -0.400 11.540 0.400 ;
        RECT  11.540 -0.400 12.520 1.170 ;
        RECT  12.520 -0.400 13.730 0.400 ;
        RECT  13.730 -0.400 14.130 0.560 ;
        RECT  14.130 -0.400 15.180 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.200 2.100 14.360 2.500 ;
        RECT  13.960 0.860 14.200 3.910 ;
        RECT  13.390 0.860 13.960 1.100 ;
        RECT  13.450 3.670 13.960 3.910 ;
        RECT  13.050 3.670 13.450 4.180 ;
        RECT  12.990 0.670 13.390 1.100 ;
        RECT  11.490 3.940 13.050 4.180 ;
        RECT  12.050 1.940 12.710 2.420 ;
        RECT  11.810 1.940 12.050 3.520 ;
        RECT  11.110 1.940 11.810 2.180 ;
        RECT  11.130 3.280 11.810 3.520 ;
        RECT  11.030 2.470 11.430 2.870 ;
        RECT  10.730 3.280 11.130 3.680 ;
        RECT  10.870 0.990 11.110 2.180 ;
        RECT  10.070 2.550 11.030 2.790 ;
        RECT  9.930 0.990 10.870 1.230 ;
        RECT  9.810 1.520 10.070 2.920 ;
        RECT  9.670 1.520 9.810 1.980 ;
        RECT  8.990 2.680 9.810 2.920 ;
        RECT  8.370 1.520 9.670 1.760 ;
        RECT  8.470 2.100 9.290 2.340 ;
        RECT  7.950 3.890 8.820 4.130 ;
        RECT  8.230 2.100 8.470 3.610 ;
        RECT  8.130 0.670 8.370 1.760 ;
        RECT  7.800 2.680 8.230 2.920 ;
        RECT  7.770 0.670 8.130 1.100 ;
        RECT  7.710 3.460 7.950 4.130 ;
        RECT  7.560 1.380 7.800 2.920 ;
        RECT  6.120 0.860 7.770 1.100 ;
        RECT  6.910 3.460 7.710 3.700 ;
        RECT  7.080 2.520 7.560 2.920 ;
        RECT  6.380 1.790 7.220 2.190 ;
        RECT  6.670 3.460 6.910 4.100 ;
        RECT  5.860 3.860 6.670 4.100 ;
        RECT  6.140 1.380 6.380 3.570 ;
        RECT  5.420 1.380 6.140 1.620 ;
        RECT  5.720 0.810 6.120 1.100 ;
        RECT  5.680 3.020 5.860 4.100 ;
        RECT  5.620 1.910 5.680 4.100 ;
        RECT  5.280 1.910 5.620 3.260 ;
        RECT  5.100 3.540 5.340 3.940 ;
        RECT  5.140 1.910 5.280 2.150 ;
        RECT  2.420 3.020 5.280 3.260 ;
        RECT  4.900 0.780 5.140 2.150 ;
        RECT  3.260 3.540 5.100 3.780 ;
        RECT  2.810 0.780 4.900 1.020 ;
        RECT  1.270 2.500 4.900 2.740 ;
        RECT  4.280 1.300 4.520 1.700 ;
        RECT  2.990 1.300 4.280 1.540 ;
        RECT  2.860 3.540 3.260 4.080 ;
        RECT  2.750 1.300 2.990 1.740 ;
        RECT  2.410 0.680 2.810 1.020 ;
        RECT  0.870 2.500 1.270 3.210 ;
        RECT  0.570 2.500 0.870 2.740 ;
        RECT  0.330 1.320 0.570 2.740 ;
        RECT  0.170 1.320 0.330 1.720 ;
    END
END JKFFXL

MACRO JKFFX4
    CLASS CORE ;
    FOREIGN JKFFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFXL ;
    SIZE 20.460 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.270 1.260 17.370 2.660 ;
        RECT  17.370 1.260 17.380 2.950 ;
        RECT  17.380 1.150 17.780 3.070 ;
        RECT  17.780 1.350 17.790 2.950 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.590 1.260 18.720 2.660 ;
        RECT  18.720 1.150 18.800 2.660 ;
        RECT  18.800 1.150 19.120 3.070 ;
        RECT  19.120 1.350 19.130 3.070 ;
        RECT  19.130 2.830 19.320 3.070 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.510 2.090 ;
        RECT  3.510 1.830 3.760 2.100 ;
        RECT  3.760 1.860 4.220 2.100 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.090 1.790 2.660 2.110 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 1.910 0.770 2.310 ;
        RECT  0.770 1.820 1.120 2.320 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.770 5.440 ;
        RECT  0.770 4.210 0.780 5.440 ;
        RECT  0.780 4.010 1.180 5.440 ;
        RECT  1.180 4.210 1.190 5.440 ;
        RECT  1.190 4.640 2.060 5.440 ;
        RECT  2.060 4.480 2.460 5.440 ;
        RECT  2.460 4.640 4.220 5.440 ;
        RECT  4.220 4.480 4.620 5.440 ;
        RECT  4.620 4.640 7.670 5.440 ;
        RECT  7.670 4.480 8.070 5.440 ;
        RECT  8.070 4.640 9.540 5.440 ;
        RECT  9.540 4.480 10.520 5.440 ;
        RECT  10.520 4.640 12.790 5.440 ;
        RECT  12.790 4.480 13.190 5.440 ;
        RECT  13.190 4.640 15.170 5.440 ;
        RECT  15.170 4.480 15.570 5.440 ;
        RECT  15.570 4.640 16.620 5.440 ;
        RECT  16.620 3.910 17.020 5.440 ;
        RECT  17.020 4.640 18.140 5.440 ;
        RECT  18.140 4.030 18.150 5.440 ;
        RECT  18.150 3.910 18.550 5.440 ;
        RECT  18.550 4.030 18.560 5.440 ;
        RECT  18.560 4.640 19.530 5.440 ;
        RECT  19.530 4.040 19.540 5.440 ;
        RECT  19.540 3.920 19.940 5.440 ;
        RECT  19.940 4.040 19.950 5.440 ;
        RECT  19.950 4.640 20.460 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.910 0.400 ;
        RECT  0.910 -0.400 1.310 0.560 ;
        RECT  1.310 -0.400 3.590 0.400 ;
        RECT  3.590 -0.400 3.990 0.560 ;
        RECT  3.990 -0.400 6.730 0.400 ;
        RECT  6.730 -0.400 7.130 0.560 ;
        RECT  7.130 -0.400 9.100 0.400 ;
        RECT  9.100 -0.400 9.110 1.060 ;
        RECT  9.110 -0.400 9.510 1.260 ;
        RECT  9.510 -0.400 9.520 1.060 ;
        RECT  9.520 -0.400 11.710 0.400 ;
        RECT  11.710 -0.400 11.720 0.740 ;
        RECT  11.720 -0.400 12.120 0.940 ;
        RECT  12.120 -0.400 12.130 0.740 ;
        RECT  12.130 -0.400 14.730 0.400 ;
        RECT  14.730 -0.400 15.130 1.040 ;
        RECT  15.130 -0.400 16.740 0.400 ;
        RECT  16.740 -0.400 16.750 0.670 ;
        RECT  16.750 -0.400 17.150 0.870 ;
        RECT  17.150 -0.400 17.160 0.670 ;
        RECT  17.160 -0.400 18.040 0.400 ;
        RECT  18.040 -0.400 18.050 0.670 ;
        RECT  18.050 -0.400 18.450 0.870 ;
        RECT  18.450 -0.400 18.460 0.670 ;
        RECT  18.460 -0.400 19.350 0.400 ;
        RECT  19.350 -0.400 19.360 0.670 ;
        RECT  19.360 -0.400 19.760 0.870 ;
        RECT  19.760 -0.400 19.770 0.670 ;
        RECT  19.770 -0.400 20.460 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  19.600 2.180 19.840 3.590 ;
        RECT  17.000 3.350 19.600 3.590 ;
        RECT  16.760 1.170 17.000 3.590 ;
        RECT  16.430 1.170 16.760 1.410 ;
        RECT  16.130 2.820 16.760 3.220 ;
        RECT  15.450 1.990 16.480 2.390 ;
        RECT  16.030 0.920 16.430 1.410 ;
        RECT  15.890 2.820 16.130 4.060 ;
        RECT  12.460 3.820 15.890 4.060 ;
        RECT  15.210 1.280 15.450 3.460 ;
        RECT  13.610 1.280 15.210 1.520 ;
        RECT  11.910 3.220 15.210 3.460 ;
        RECT  14.630 2.490 14.790 2.730 ;
        RECT  14.390 1.760 14.630 2.730 ;
        RECT  13.120 1.760 14.390 2.000 ;
        RECT  13.950 2.240 14.110 2.480 ;
        RECT  13.710 2.240 13.950 2.870 ;
        RECT  11.160 2.630 13.710 2.870 ;
        RECT  13.210 1.030 13.610 1.520 ;
        RECT  11.430 1.280 13.210 1.520 ;
        RECT  12.880 1.760 13.120 2.080 ;
        RECT  10.490 1.840 12.880 2.080 ;
        RECT  12.220 3.820 12.460 4.180 ;
        RECT  7.390 3.940 12.220 4.180 ;
        RECT  11.510 3.220 11.910 3.640 ;
        RECT  11.190 1.020 11.430 1.520 ;
        RECT  10.730 1.020 11.190 1.260 ;
        RECT  10.920 2.630 11.160 3.590 ;
        RECT  6.870 3.350 10.920 3.590 ;
        RECT  10.330 0.860 10.730 1.260 ;
        RECT  10.480 1.630 10.490 2.080 ;
        RECT  10.320 1.540 10.480 2.080 ;
        RECT  10.080 1.540 10.320 2.980 ;
        RECT  8.750 1.540 10.080 1.780 ;
        RECT  9.440 2.740 10.080 2.980 ;
        RECT  9.310 2.060 9.710 2.460 ;
        RECT  8.640 2.220 9.310 2.460 ;
        RECT  8.510 0.860 8.750 1.780 ;
        RECT  8.480 2.220 8.640 3.060 ;
        RECT  8.350 0.860 8.510 1.290 ;
        RECT  8.240 2.210 8.480 3.060 ;
        RECT  6.450 0.860 8.350 1.100 ;
        RECT  8.070 2.210 8.240 2.580 ;
        RECT  7.830 1.380 8.070 2.580 ;
        RECT  7.610 1.380 7.830 1.620 ;
        RECT  7.450 2.340 7.830 2.580 ;
        RECT  7.050 2.330 7.450 2.730 ;
        RECT  7.150 3.940 7.390 4.360 ;
        RECT  7.080 1.610 7.320 2.020 ;
        RECT  5.300 4.120 7.150 4.360 ;
        RECT  6.350 1.620 7.080 2.020 ;
        RECT  6.630 3.350 6.870 3.840 ;
        RECT  5.830 3.600 6.630 3.840 ;
        RECT  6.210 0.680 6.450 1.100 ;
        RECT  6.110 1.400 6.350 3.330 ;
        RECT  5.840 0.680 6.210 0.920 ;
        RECT  5.840 1.400 6.110 1.640 ;
        RECT  5.600 1.240 5.840 1.640 ;
        RECT  5.660 2.900 5.830 3.840 ;
        RECT  5.590 1.920 5.660 3.840 ;
        RECT  5.260 1.920 5.590 3.140 ;
        RECT  2.930 3.420 5.310 3.660 ;
        RECT  5.060 3.940 5.300 4.360 ;
        RECT  2.580 2.900 5.260 3.140 ;
        RECT  3.580 3.940 5.060 4.180 ;
        RECT  2.060 2.380 4.940 2.620 ;
        RECT  2.840 1.280 4.700 1.520 ;
        RECT  3.180 3.940 3.580 4.370 ;
        RECT  1.460 3.940 3.180 4.180 ;
        RECT  2.340 2.900 2.580 3.550 ;
        RECT  1.820 1.280 2.500 1.520 ;
        RECT  0.580 3.310 2.340 3.550 ;
        RECT  1.820 2.380 2.060 3.010 ;
        RECT  1.580 1.280 1.820 3.010 ;
        RECT  0.570 3.130 0.580 3.550 ;
        RECT  0.400 2.850 0.570 3.550 ;
        RECT  0.400 1.200 0.490 1.600 ;
        RECT  0.160 1.200 0.400 3.550 ;
    END
END JKFFX4

MACRO JKFFX2
    CLASS CORE ;
    FOREIGN JKFFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFXL ;
    SIZE 17.820 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.000 1.170 15.300 1.570 ;
        RECT  15.300 1.170 15.400 3.410 ;
        RECT  15.400 1.330 15.540 3.410 ;
        RECT  15.540 2.950 15.640 3.410 ;
        RECT  15.640 2.960 15.790 3.410 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.700 2.390 16.710 2.650 ;
        RECT  16.440 1.070 16.710 1.470 ;
        RECT  16.710 1.070 16.950 3.340 ;
        RECT  16.950 2.390 16.960 2.650 ;
        RECT  16.950 3.100 17.030 3.340 ;
        RECT  17.030 3.100 17.430 3.500 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.410 1.820 3.760 2.210 ;
        RECT  3.760 1.960 3.940 2.200 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.520 0.700 0.770 1.100 ;
        RECT  0.770 0.700 0.860 1.510 ;
        RECT  0.860 0.700 0.920 1.530 ;
        RECT  0.920 0.860 1.010 1.530 ;
        RECT  1.010 1.270 1.120 1.530 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.800 1.870 2.090 ;
        RECT  1.870 1.800 2.270 2.200 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.370 5.440 ;
        RECT  0.370 3.830 0.380 5.440 ;
        RECT  0.380 3.630 0.780 5.440 ;
        RECT  0.780 3.830 0.790 5.440 ;
        RECT  0.790 4.640 1.540 5.440 ;
        RECT  1.540 3.470 1.550 5.440 ;
        RECT  1.550 3.270 1.950 5.440 ;
        RECT  1.950 3.470 1.960 5.440 ;
        RECT  1.960 4.640 4.070 5.440 ;
        RECT  4.070 4.160 4.080 5.440 ;
        RECT  4.080 4.040 4.480 5.440 ;
        RECT  4.480 4.160 4.490 5.440 ;
        RECT  4.490 4.640 7.150 5.440 ;
        RECT  7.150 4.310 7.160 5.440 ;
        RECT  7.160 4.110 7.560 5.440 ;
        RECT  7.560 4.310 7.570 5.440 ;
        RECT  7.570 4.640 9.590 5.440 ;
        RECT  9.590 4.200 9.600 5.440 ;
        RECT  9.600 4.000 10.000 5.440 ;
        RECT  10.000 4.200 10.010 5.440 ;
        RECT  10.010 4.640 12.110 5.440 ;
        RECT  12.110 4.120 12.120 5.440 ;
        RECT  12.120 3.920 12.520 5.440 ;
        RECT  12.520 4.120 12.530 5.440 ;
        RECT  12.530 4.640 13.940 5.440 ;
        RECT  13.940 4.480 14.340 5.440 ;
        RECT  14.340 4.640 16.200 5.440 ;
        RECT  16.200 4.350 16.210 5.440 ;
        RECT  16.210 4.230 16.610 5.440 ;
        RECT  16.610 4.350 16.620 5.440 ;
        RECT  16.620 4.640 17.820 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.500 0.400 ;
        RECT  1.500 -0.400 1.900 0.560 ;
        RECT  1.900 -0.400 6.450 0.400 ;
        RECT  6.450 -0.400 7.430 0.560 ;
        RECT  7.430 -0.400 8.700 0.400 ;
        RECT  8.700 -0.400 8.710 0.800 ;
        RECT  8.710 -0.400 9.110 1.000 ;
        RECT  9.110 -0.400 9.120 0.800 ;
        RECT  9.120 -0.400 11.170 0.400 ;
        RECT  11.170 -0.400 11.570 0.560 ;
        RECT  11.570 -0.400 13.320 0.400 ;
        RECT  13.320 -0.400 13.720 0.560 ;
        RECT  13.720 -0.400 15.710 0.400 ;
        RECT  15.710 -0.400 15.720 0.860 ;
        RECT  15.720 -0.400 16.120 1.060 ;
        RECT  16.120 -0.400 16.130 0.860 ;
        RECT  16.130 -0.400 17.820 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.100 1.780 16.340 3.930 ;
        RECT  15.940 1.780 16.100 2.180 ;
        RECT  15.010 3.690 16.100 3.930 ;
        RECT  14.850 1.860 15.010 3.930 ;
        RECT  14.770 1.860 14.850 4.170 ;
        RECT  14.520 1.860 14.770 2.100 ;
        RECT  14.590 3.060 14.770 4.170 ;
        RECT  13.650 3.930 14.590 4.170 ;
        RECT  14.280 1.010 14.520 2.100 ;
        RECT  13.740 2.380 14.490 2.780 ;
        RECT  14.120 1.010 14.280 1.410 ;
        RECT  13.500 0.900 13.740 3.500 ;
        RECT  13.330 3.930 13.650 4.350 ;
        RECT  12.380 0.900 13.500 1.140 ;
        RECT  13.010 3.260 13.500 3.500 ;
        RECT  13.250 3.950 13.330 4.350 ;
        RECT  12.980 1.440 13.220 2.920 ;
        RECT  12.600 3.260 13.010 3.520 ;
        RECT  10.070 1.440 12.980 1.680 ;
        RECT  12.820 2.680 12.980 2.920 ;
        RECT  11.220 1.960 12.700 2.200 ;
        RECT  11.260 3.280 12.600 3.520 ;
        RECT  11.980 0.900 12.380 1.160 ;
        RECT  10.310 0.900 11.980 1.140 ;
        RECT  10.860 3.280 11.260 3.680 ;
        RECT  11.220 2.480 11.230 2.880 ;
        RECT  10.980 1.960 11.220 2.880 ;
        RECT  10.830 2.480 10.980 2.880 ;
        RECT  10.570 2.640 10.830 2.880 ;
        RECT  10.330 2.640 10.570 3.710 ;
        RECT  9.320 3.470 10.330 3.710 ;
        RECT  9.910 0.740 10.310 1.140 ;
        RECT  9.920 1.420 10.070 1.830 ;
        RECT  9.680 1.420 9.920 3.190 ;
        RECT  9.670 1.420 9.680 1.830 ;
        RECT  8.800 2.950 9.680 3.190 ;
        RECT  8.430 1.420 9.670 1.670 ;
        RECT  8.930 3.470 9.320 3.980 ;
        RECT  8.500 1.950 9.290 2.190 ;
        RECT  8.920 3.550 8.930 3.980 ;
        RECT  6.870 3.550 8.920 3.790 ;
        RECT  8.440 1.950 8.500 3.070 ;
        RECT  8.260 1.950 8.440 3.310 ;
        RECT  8.190 0.670 8.430 1.670 ;
        RECT  8.040 2.830 8.260 3.310 ;
        RECT  7.830 0.670 8.190 1.100 ;
        RECT  7.810 2.830 8.040 3.070 ;
        RECT  6.180 0.860 7.830 1.100 ;
        RECT  7.570 1.380 7.810 3.070 ;
        RECT  7.020 2.670 7.570 3.070 ;
        RECT  6.320 1.950 7.290 2.350 ;
        RECT  6.630 3.550 6.870 4.270 ;
        RECT  5.800 4.030 6.630 4.270 ;
        RECT  6.080 1.380 6.320 3.720 ;
        RECT  5.780 0.810 6.180 1.100 ;
        RECT  5.480 1.380 6.080 1.620 ;
        RECT  5.580 3.000 5.800 4.270 ;
        RECT  5.560 1.910 5.580 4.270 ;
        RECT  5.190 1.910 5.560 3.240 ;
        RECT  5.040 3.520 5.280 3.920 ;
        RECT  5.180 1.910 5.190 2.310 ;
        RECT  2.270 3.000 5.190 3.240 ;
        RECT  5.140 1.910 5.180 2.150 ;
        RECT  4.900 0.780 5.140 2.150 ;
        RECT  3.220 3.520 5.040 3.760 ;
        RECT  2.710 0.780 4.900 1.020 ;
        RECT  1.010 2.480 4.840 2.720 ;
        RECT  4.220 1.300 4.460 1.700 ;
        RECT  2.810 1.300 4.220 1.540 ;
        RECT  2.820 3.520 3.220 4.060 ;
        RECT  2.570 1.300 2.810 1.830 ;
        RECT  2.310 0.680 2.710 1.020 ;
        RECT  0.610 2.480 1.010 3.160 ;
        RECT  0.410 2.480 0.610 2.720 ;
        RECT  0.410 1.380 0.490 1.780 ;
        RECT  0.170 1.380 0.410 2.720 ;
    END
END JKFFX2

MACRO JKFFX1
    CLASS CORE ;
    FOREIGN JKFFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ JKFFXL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.920 3.970 13.080 4.370 ;
        RECT  12.910 0.690 13.310 1.100 ;
        RECT  13.080 3.530 13.320 4.370 ;
        RECT  13.320 3.530 13.400 3.770 ;
        RECT  13.400 3.510 13.420 3.770 ;
        RECT  13.420 3.500 13.660 3.770 ;
        RECT  13.660 3.500 13.820 3.740 ;
        RECT  13.310 0.860 13.820 1.100 ;
        RECT  13.820 0.860 14.060 3.740 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.580 1.780 14.590 3.080 ;
        RECT  14.590 1.390 14.990 3.240 ;
        RECT  14.990 1.780 15.000 3.080 ;
        END
    END Q
    PIN K
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.410 1.820 3.760 2.210 ;
        RECT  3.760 1.960 3.940 2.200 ;
        END
    END K
    PIN J
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.570 3.500 0.850 3.900 ;
        RECT  0.850 3.490 1.120 3.910 ;
        END
    END J
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.800 1.840 2.090 ;
        RECT  1.840 1.800 2.240 2.200 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.740 5.440 ;
        RECT  1.740 3.920 1.750 5.440 ;
        RECT  1.750 3.720 2.150 5.440 ;
        RECT  2.150 3.920 2.160 5.440 ;
        RECT  2.160 4.640 4.130 5.440 ;
        RECT  4.130 4.160 4.140 5.440 ;
        RECT  4.140 4.040 4.540 5.440 ;
        RECT  4.540 4.160 4.550 5.440 ;
        RECT  4.550 4.640 7.190 5.440 ;
        RECT  7.190 3.980 7.430 5.440 ;
        RECT  7.430 4.640 9.280 5.440 ;
        RECT  9.280 3.930 9.290 5.440 ;
        RECT  9.290 3.730 9.690 5.440 ;
        RECT  9.690 3.930 9.700 5.440 ;
        RECT  9.700 4.640 12.120 5.440 ;
        RECT  12.120 4.480 12.520 5.440 ;
        RECT  12.520 4.640 13.780 5.440 ;
        RECT  13.780 4.480 14.180 5.440 ;
        RECT  14.180 4.640 15.180 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.500 0.400 ;
        RECT  1.500 -0.400 1.900 0.560 ;
        RECT  1.900 -0.400 6.450 0.400 ;
        RECT  6.450 -0.400 7.430 0.560 ;
        RECT  7.430 -0.400 8.700 0.400 ;
        RECT  8.700 -0.400 8.710 1.110 ;
        RECT  8.710 -0.400 9.110 1.310 ;
        RECT  9.110 -0.400 9.120 1.110 ;
        RECT  9.120 -0.400 11.540 0.400 ;
        RECT  11.540 -0.400 12.520 1.170 ;
        RECT  12.520 -0.400 13.790 0.400 ;
        RECT  13.790 -0.400 14.190 0.560 ;
        RECT  14.190 -0.400 15.180 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  13.380 2.090 13.540 2.490 ;
        RECT  13.380 1.390 13.390 1.790 ;
        RECT  13.140 1.390 13.380 3.210 ;
        RECT  12.990 1.390 13.140 1.790 ;
        RECT  12.920 2.810 13.140 3.210 ;
        RECT  12.570 2.970 12.920 3.210 ;
        RECT  12.050 2.020 12.710 2.420 ;
        RECT  12.330 2.970 12.570 4.050 ;
        RECT  11.490 3.810 12.330 4.050 ;
        RECT  11.810 1.860 12.050 3.300 ;
        RECT  11.110 1.860 11.810 2.100 ;
        RECT  11.130 3.060 11.810 3.300 ;
        RECT  11.030 2.380 11.430 2.780 ;
        RECT  10.730 3.060 11.130 3.680 ;
        RECT  10.870 1.070 11.110 2.100 ;
        RECT  10.070 2.460 11.030 2.700 ;
        RECT  10.330 1.070 10.870 1.310 ;
        RECT  9.930 0.910 10.330 1.310 ;
        RECT  9.910 1.730 10.070 2.700 ;
        RECT  9.670 1.730 9.910 3.160 ;
        RECT  8.430 1.730 9.670 1.970 ;
        RECT  8.990 2.920 9.670 3.160 ;
        RECT  8.470 2.250 9.290 2.490 ;
        RECT  7.950 3.890 8.820 4.130 ;
        RECT  8.230 2.250 8.470 3.570 ;
        RECT  8.180 0.670 8.430 1.970 ;
        RECT  7.860 2.680 8.230 2.920 ;
        RECT  7.830 0.670 8.180 1.100 ;
        RECT  7.710 3.460 7.950 4.130 ;
        RECT  7.620 1.380 7.860 2.920 ;
        RECT  6.180 0.860 7.830 1.100 ;
        RECT  6.910 3.460 7.710 3.700 ;
        RECT  7.080 2.520 7.620 2.920 ;
        RECT  6.380 1.790 7.290 2.190 ;
        RECT  6.670 3.460 6.910 4.100 ;
        RECT  5.860 3.860 6.670 4.100 ;
        RECT  6.140 1.380 6.380 3.570 ;
        RECT  5.780 0.810 6.180 1.100 ;
        RECT  5.480 1.380 6.140 1.620 ;
        RECT  5.620 3.000 5.860 4.100 ;
        RECT  5.580 3.000 5.620 3.240 ;
        RECT  5.180 1.910 5.580 3.240 ;
        RECT  5.100 3.520 5.340 3.920 ;
        RECT  5.140 1.910 5.180 2.150 ;
        RECT  2.330 3.000 5.180 3.240 ;
        RECT  4.900 0.780 5.140 2.150 ;
        RECT  3.200 3.520 5.100 3.760 ;
        RECT  2.810 0.780 4.900 1.020 ;
        RECT  1.270 2.480 4.840 2.720 ;
        RECT  4.220 1.300 4.460 1.700 ;
        RECT  2.810 1.300 4.220 1.540 ;
        RECT  2.800 3.520 3.200 4.060 ;
        RECT  2.410 0.680 2.810 1.020 ;
        RECT  2.570 1.300 2.810 1.740 ;
        RECT  0.870 2.480 1.270 3.210 ;
        RECT  0.570 2.480 0.870 2.720 ;
        RECT  0.330 1.320 0.570 2.720 ;
        RECT  0.170 1.320 0.330 1.720 ;
    END
END JKFFX1

MACRO INVXL
    CLASS CORE ;
    FOREIGN INVXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 0.870 3.210 ;
        RECT  0.870 2.920 1.070 3.210 ;
        RECT  1.070 1.380 1.110 3.210 ;
        RECT  1.110 1.380 1.310 3.240 ;
        RECT  1.310 2.840 1.350 3.240 ;
        RECT  1.310 1.380 1.470 1.780 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.270 0.210 1.530 ;
        RECT  0.210 1.270 0.450 2.440 ;
        RECT  0.450 1.270 0.460 1.530 ;
        RECT  0.450 1.830 0.680 2.440 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 3.730 0.180 5.440 ;
        RECT  0.180 3.530 0.580 5.440 ;
        RECT  0.580 3.730 0.590 5.440 ;
        RECT  0.590 4.640 1.980 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.070 0.400 ;
        RECT  1.070 -0.400 1.470 0.560 ;
        RECT  1.470 -0.400 1.980 0.400 ;
        END
    END GND
END INVXL

MACRO INVX8
    CLASS CORE ;
    FOREIGN INVX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ INVXL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.760 2.930 1.520 3.410 ;
        RECT  0.750 1.250 1.520 1.730 ;
        RECT  1.520 1.250 3.100 3.410 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.300 2.180 0.850 2.580 ;
        RECT  0.850 2.180 0.860 2.640 ;
        RECT  0.860 2.180 1.120 2.650 ;
        RECT  1.120 2.180 1.280 2.580 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.180 5.440 ;
        RECT  0.180 4.120 0.190 5.440 ;
        RECT  0.190 3.920 0.590 5.440 ;
        RECT  0.590 4.120 0.600 5.440 ;
        RECT  0.600 4.640 1.660 5.440 ;
        RECT  1.660 4.120 1.670 5.440 ;
        RECT  1.670 3.920 2.070 5.440 ;
        RECT  2.070 4.120 2.080 5.440 ;
        RECT  2.080 4.640 3.020 5.440 ;
        RECT  3.020 4.220 3.030 5.440 ;
        RECT  3.030 4.020 3.430 5.440 ;
        RECT  3.430 4.220 3.440 5.440 ;
        RECT  3.440 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 0.780 ;
        RECT  0.170 -0.400 0.570 0.980 ;
        RECT  0.570 -0.400 0.580 0.780 ;
        RECT  0.580 -0.400 1.490 0.400 ;
        RECT  1.490 -0.400 1.500 0.780 ;
        RECT  1.500 -0.400 1.900 0.980 ;
        RECT  1.900 -0.400 1.910 0.780 ;
        RECT  1.910 -0.400 2.910 0.400 ;
        RECT  2.910 -0.400 3.310 0.560 ;
        RECT  3.310 -0.400 4.620 0.400 ;
        END
    END GND
END INVX8

MACRO INVX4
    CLASS CORE ;
    FOREIGN INVX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ INVXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.310 1.160 1.330 1.560 ;
        RECT  1.330 1.140 1.430 1.560 ;
        RECT  1.430 1.140 1.440 3.220 ;
        RECT  1.440 1.140 1.790 3.250 ;
        RECT  1.790 1.820 1.840 3.250 ;
        RECT  1.840 1.820 1.870 3.220 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.210 2.650 ;
        RECT  0.210 2.060 0.460 2.650 ;
        RECT  0.460 2.060 0.760 2.470 ;
        RECT  0.760 2.070 1.160 2.470 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.740 5.440 ;
        RECT  0.740 4.000 0.750 5.440 ;
        RECT  0.750 3.800 1.150 5.440 ;
        RECT  1.150 4.000 1.160 5.440 ;
        RECT  1.160 4.640 2.060 5.440 ;
        RECT  2.060 4.210 2.070 5.440 ;
        RECT  2.070 4.010 2.470 5.440 ;
        RECT  2.470 4.210 2.480 5.440 ;
        RECT  2.480 4.640 2.640 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.540 0.400 ;
        RECT  0.540 -0.400 0.550 1.310 ;
        RECT  0.550 -0.400 0.950 1.510 ;
        RECT  0.950 -0.400 0.960 1.310 ;
        RECT  0.960 -0.400 2.060 0.400 ;
        RECT  2.060 -0.400 2.070 1.070 ;
        RECT  2.070 -0.400 2.470 1.560 ;
        RECT  2.470 -0.400 2.480 1.070 ;
        RECT  2.480 -0.400 2.640 0.400 ;
        END
    END GND
END INVX4

MACRO INVX3
    CLASS CORE ;
    FOREIGN INVX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ INVXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.770 2.940 0.870 3.780 ;
        RECT  0.870 2.750 0.980 3.780 ;
        RECT  0.980 2.740 1.140 3.780 ;
        RECT  0.980 1.110 1.140 1.760 ;
        RECT  1.140 1.110 1.210 3.780 ;
        RECT  1.210 1.110 1.380 3.720 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.220 2.650 ;
        RECT  0.220 2.200 0.230 2.650 ;
        RECT  0.230 2.040 0.460 2.650 ;
        RECT  0.460 2.040 0.900 2.440 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 1.710 5.440 ;
        RECT  1.710 3.480 1.720 5.440 ;
        RECT  1.720 3.000 2.120 5.440 ;
        RECT  2.120 3.480 2.130 5.440 ;
        RECT  2.130 4.640 2.640 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 1.710 0.400 ;
        RECT  1.710 -0.400 1.720 1.270 ;
        RECT  1.720 -0.400 2.120 1.470 ;
        RECT  2.120 -0.400 2.130 1.270 ;
        RECT  2.130 -0.400 2.640 0.400 ;
        END
    END GND
END INVX3

MACRO INVX2
    CLASS CORE ;
    FOREIGN INVX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ INVXL ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.190 1.390 1.350 1.790 ;
        RECT  0.780 3.100 1.530 3.520 ;
        RECT  1.520 2.390 1.530 2.650 ;
        RECT  1.350 1.390 1.530 1.820 ;
        RECT  1.530 1.390 1.590 3.520 ;
        RECT  1.590 1.580 1.770 3.520 ;
        RECT  1.770 3.070 1.780 3.520 ;
        RECT  1.770 2.390 1.780 2.650 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.460 2.510 ;
        RECT  0.460 2.100 0.550 2.510 ;
        RECT  0.550 2.110 1.160 2.510 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.060 5.440 ;
        RECT  1.060 4.480 1.460 5.440 ;
        RECT  1.460 4.640 1.980 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.180 0.400 ;
        RECT  1.180 -0.400 1.190 0.870 ;
        RECT  1.190 -0.400 1.590 1.070 ;
        RECT  1.590 -0.400 1.600 0.870 ;
        RECT  1.600 -0.400 1.980 0.400 ;
        END
    END GND
END INVX2

MACRO INVX20
    CLASS CORE ;
    FOREIGN INVX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ INVXL ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  5.720 2.840 6.230 3.820 ;
        RECT  6.230 2.840 6.930 3.520 ;
        RECT  6.930 2.840 7.670 3.820 ;
        RECT  7.670 2.840 8.810 3.520 ;
        RECT  8.810 2.840 9.570 3.820 ;
        RECT  9.570 2.840 9.850 3.520 ;
        RECT  9.850 2.510 10.110 3.520 ;
        RECT  5.580 1.200 10.110 1.880 ;
        RECT  10.110 1.200 11.670 3.840 ;
        RECT  11.670 2.510 11.930 3.820 ;
        RECT  11.930 2.840 12.290 3.820 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.060 0.460 2.650 ;
        RECT  0.460 2.060 0.750 2.480 ;
        RECT  0.750 2.070 0.960 2.470 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.600 0.560 5.440 ;
        RECT  0.560 4.640 1.500 5.440 ;
        RECT  1.500 4.130 1.900 5.440 ;
        RECT  1.900 4.640 3.090 5.440 ;
        RECT  3.090 4.130 3.490 5.440 ;
        RECT  3.490 4.640 4.710 5.440 ;
        RECT  4.710 3.000 5.110 5.440 ;
        RECT  5.110 4.480 5.450 5.440 ;
        RECT  5.450 4.640 6.510 5.440 ;
        RECT  6.510 4.360 6.520 5.440 ;
        RECT  6.520 4.160 6.920 5.440 ;
        RECT  6.920 4.360 6.930 5.440 ;
        RECT  6.930 4.640 8.060 5.440 ;
        RECT  8.060 4.360 8.070 5.440 ;
        RECT  8.070 4.160 8.470 5.440 ;
        RECT  8.470 4.360 8.480 5.440 ;
        RECT  8.480 4.640 9.610 5.440 ;
        RECT  9.610 4.360 9.620 5.440 ;
        RECT  9.620 4.160 10.020 5.440 ;
        RECT  10.020 4.360 10.030 5.440 ;
        RECT  10.030 4.640 11.150 5.440 ;
        RECT  11.150 4.350 11.160 5.440 ;
        RECT  11.160 4.150 11.560 5.440 ;
        RECT  11.560 4.350 11.570 5.440 ;
        RECT  11.570 4.640 12.540 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 1.300 ;
        RECT  0.170 -0.400 0.570 1.500 ;
        RECT  0.570 -0.400 0.580 1.300 ;
        RECT  0.580 -0.400 1.690 0.400 ;
        RECT  1.690 -0.400 1.700 0.850 ;
        RECT  1.700 -0.400 2.100 1.050 ;
        RECT  2.100 -0.400 2.110 0.850 ;
        RECT  2.110 -0.400 3.030 0.400 ;
        RECT  3.030 -0.400 3.040 0.850 ;
        RECT  3.040 -0.400 3.440 1.050 ;
        RECT  3.440 -0.400 3.450 0.850 ;
        RECT  3.450 -0.400 4.680 0.400 ;
        RECT  4.680 -0.400 5.080 1.780 ;
        RECT  5.080 -0.400 5.380 0.560 ;
        RECT  5.380 -0.400 6.380 0.400 ;
        RECT  6.380 -0.400 6.390 0.810 ;
        RECT  6.390 -0.400 6.790 0.930 ;
        RECT  6.790 -0.400 6.800 0.810 ;
        RECT  6.800 -0.400 7.720 0.400 ;
        RECT  7.720 -0.400 7.730 0.780 ;
        RECT  7.730 -0.400 8.130 0.900 ;
        RECT  8.130 -0.400 8.140 0.780 ;
        RECT  8.140 -0.400 9.060 0.400 ;
        RECT  9.060 -0.400 9.070 0.780 ;
        RECT  9.070 -0.400 9.470 0.900 ;
        RECT  9.470 -0.400 9.480 0.780 ;
        RECT  9.480 -0.400 10.400 0.400 ;
        RECT  10.400 -0.400 10.410 0.780 ;
        RECT  10.410 -0.400 10.810 0.900 ;
        RECT  10.810 -0.400 10.820 0.780 ;
        RECT  10.820 -0.400 12.540 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.530 2.160 9.610 2.560 ;
        RECT  4.140 2.210 5.530 2.510 ;
        RECT  4.050 1.490 4.140 3.290 ;
        RECT  3.840 1.390 4.050 3.290 ;
        RECT  2.370 1.390 3.840 1.790 ;
        RECT  3.740 2.840 3.840 3.290 ;
        RECT  2.670 2.840 3.740 3.140 ;
        RECT  1.500 2.070 3.600 2.470 ;
        RECT  2.270 2.840 2.670 3.820 ;
        RECT  1.260 1.390 1.500 2.990 ;
        RECT  0.970 1.390 1.260 1.790 ;
        RECT  1.220 2.750 1.260 2.990 ;
        RECT  0.820 2.750 1.220 3.150 ;
    END
END INVX20

MACRO INVX1
    CLASS CORE ;
    FOREIGN INVX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ INVXL ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 1.040 3.210 ;
        RECT  1.040 1.280 1.280 3.240 ;
        RECT  1.280 2.840 1.440 3.240 ;
        RECT  1.280 1.280 1.440 1.680 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.430 2.090 ;
        RECT  0.430 1.830 0.460 2.580 ;
        RECT  0.460 1.850 0.670 2.580 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.200 5.440 ;
        RECT  0.200 3.690 0.210 5.440 ;
        RECT  0.210 3.490 0.610 5.440 ;
        RECT  0.610 3.690 0.620 5.440 ;
        RECT  0.620 4.640 1.980 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.980 0.400 ;
        END
    END GND
END INVX1

MACRO INVX16
    CLASS CORE ;
    FOREIGN INVX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ INVXL ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  5.520 1.200 6.950 1.880 ;
        RECT  6.950 0.840 7.350 1.880 ;
        RECT  5.290 2.840 7.870 3.840 ;
        RECT  7.870 2.520 8.130 3.840 ;
        RECT  7.350 1.200 8.130 1.880 ;
        RECT  8.130 1.200 8.490 3.840 ;
        RECT  8.490 0.840 8.890 3.840 ;
        RECT  8.890 1.200 9.690 3.840 ;
        RECT  9.690 1.200 10.300 1.930 ;
        RECT  9.690 2.520 10.310 3.840 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.720 2.070 0.860 2.470 ;
        RECT  0.860 2.070 1.120 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.190 5.440 ;
        RECT  0.190 3.130 0.200 5.440 ;
        RECT  0.200 2.930 0.600 5.440 ;
        RECT  0.600 3.130 0.610 5.440 ;
        RECT  0.610 4.640 1.550 5.440 ;
        RECT  1.550 4.000 1.950 5.440 ;
        RECT  1.950 4.640 2.980 5.440 ;
        RECT  2.980 4.100 2.990 5.440 ;
        RECT  2.990 3.620 3.390 5.440 ;
        RECT  3.390 4.100 3.400 5.440 ;
        RECT  3.400 4.640 4.530 5.440 ;
        RECT  4.530 4.100 4.540 5.440 ;
        RECT  4.540 3.620 4.940 5.440 ;
        RECT  4.940 4.100 4.950 5.440 ;
        RECT  4.950 4.640 6.110 5.440 ;
        RECT  6.110 4.360 6.120 5.440 ;
        RECT  6.120 4.160 6.520 5.440 ;
        RECT  6.520 4.360 6.530 5.440 ;
        RECT  6.530 4.640 7.660 5.440 ;
        RECT  7.660 4.360 7.670 5.440 ;
        RECT  7.670 4.160 8.070 5.440 ;
        RECT  8.070 4.360 8.080 5.440 ;
        RECT  8.080 4.640 9.200 5.440 ;
        RECT  9.200 4.360 9.210 5.440 ;
        RECT  9.210 4.160 9.610 5.440 ;
        RECT  9.610 4.360 9.620 5.440 ;
        RECT  9.620 4.640 10.560 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.740 0.400 ;
        RECT  1.740 -0.400 1.750 0.850 ;
        RECT  1.750 -0.400 2.150 1.050 ;
        RECT  2.150 -0.400 2.160 0.850 ;
        RECT  2.160 -0.400 3.120 0.400 ;
        RECT  3.120 -0.400 3.130 0.850 ;
        RECT  3.130 -0.400 3.530 1.050 ;
        RECT  3.530 -0.400 3.540 0.850 ;
        RECT  3.540 -0.400 4.790 0.400 ;
        RECT  4.790 -0.400 4.800 1.250 ;
        RECT  4.800 -0.400 5.200 1.450 ;
        RECT  5.200 -0.400 5.210 1.250 ;
        RECT  5.210 -0.400 6.140 0.400 ;
        RECT  6.140 -0.400 6.150 0.730 ;
        RECT  6.150 -0.400 6.550 0.930 ;
        RECT  6.550 -0.400 6.560 0.730 ;
        RECT  6.560 -0.400 7.680 0.400 ;
        RECT  7.680 -0.400 7.690 0.730 ;
        RECT  7.690 -0.400 8.090 0.930 ;
        RECT  8.090 -0.400 8.100 0.730 ;
        RECT  8.100 -0.400 9.210 0.400 ;
        RECT  9.210 -0.400 9.220 0.730 ;
        RECT  9.220 -0.400 9.620 0.930 ;
        RECT  9.620 -0.400 9.630 0.730 ;
        RECT  9.630 -0.400 10.560 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.460 2.160 7.630 2.560 ;
        RECT  4.140 1.390 4.460 3.300 ;
        RECT  4.060 1.390 4.140 3.840 ;
        RECT  2.460 1.390 4.060 1.790 ;
        RECT  3.740 2.880 4.060 3.840 ;
        RECT  2.210 2.070 3.770 2.470 ;
        RECT  2.270 2.890 3.740 3.290 ;
        RECT  1.880 2.070 2.210 2.310 ;
        RECT  1.640 1.550 1.880 3.170 ;
        RECT  1.500 1.550 1.640 1.790 ;
        RECT  1.360 2.930 1.640 3.170 ;
        RECT  1.100 1.390 1.500 1.790 ;
        RECT  0.960 2.930 1.360 3.330 ;
    END
END INVX16

MACRO INVX12
    CLASS CORE ;
    FOREIGN INVX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ INVXL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.170 2.860 6.150 3.540 ;
        RECT  4.150 1.200 6.150 1.880 ;
        RECT  6.150 1.200 7.510 3.840 ;
        RECT  7.510 1.520 7.710 3.840 ;
        RECT  7.710 1.520 7.720 1.960 ;
        RECT  7.710 3.050 7.770 3.640 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.080 0.780 2.480 ;
        RECT  0.780 1.840 0.860 2.480 ;
        RECT  0.860 1.830 1.020 2.480 ;
        RECT  1.020 1.830 1.120 2.090 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.880 5.440 ;
        RECT  0.880 4.130 1.280 5.440 ;
        RECT  1.280 4.640 2.340 5.440 ;
        RECT  2.340 4.480 2.740 5.440 ;
        RECT  2.740 4.640 3.620 5.440 ;
        RECT  3.620 4.480 4.020 5.440 ;
        RECT  4.020 4.640 5.100 5.440 ;
        RECT  5.100 4.360 5.110 5.440 ;
        RECT  5.110 4.160 5.510 5.440 ;
        RECT  5.510 4.360 5.520 5.440 ;
        RECT  5.520 4.640 6.660 5.440 ;
        RECT  6.660 4.360 6.670 5.440 ;
        RECT  6.670 4.160 7.070 5.440 ;
        RECT  7.070 4.360 7.080 5.440 ;
        RECT  7.080 4.640 8.020 5.440 ;
        RECT  8.020 4.160 8.420 5.440 ;
        RECT  8.420 4.640 8.580 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.910 0.400 ;
        RECT  0.910 -0.400 1.310 1.030 ;
        RECT  1.310 -0.400 2.290 0.400 ;
        RECT  2.290 -0.400 2.690 0.560 ;
        RECT  2.690 -0.400 3.620 0.400 ;
        RECT  3.620 -0.400 4.020 0.560 ;
        RECT  4.020 -0.400 4.950 0.400 ;
        RECT  4.950 -0.400 4.960 0.730 ;
        RECT  4.960 -0.400 5.360 0.930 ;
        RECT  5.360 -0.400 5.370 0.730 ;
        RECT  5.370 -0.400 6.290 0.400 ;
        RECT  6.290 -0.400 6.300 0.730 ;
        RECT  6.300 -0.400 6.700 0.930 ;
        RECT  6.700 -0.400 6.710 0.730 ;
        RECT  6.710 -0.400 8.580 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.280 2.160 5.820 2.560 ;
        RECT  3.430 2.210 4.280 2.510 ;
        RECT  3.430 2.890 3.440 3.290 ;
        RECT  3.420 2.210 3.430 3.290 ;
        RECT  3.340 1.390 3.420 3.290 ;
        RECT  3.130 1.390 3.340 3.570 ;
        RECT  3.120 1.390 3.130 2.510 ;
        RECT  3.040 2.890 3.130 3.570 ;
        RECT  3.020 1.390 3.120 1.800 ;
        RECT  2.080 3.270 3.040 3.570 ;
        RECT  2.020 1.500 3.020 1.800 ;
        RECT  1.990 2.070 2.860 2.470 ;
        RECT  1.730 3.270 2.080 3.680 ;
        RECT  1.670 1.390 2.020 1.800 ;
        RECT  1.880 2.070 1.990 3.000 ;
        RECT  1.750 2.150 1.880 3.000 ;
        RECT  0.560 2.760 1.750 3.000 ;
        RECT  1.680 3.280 1.730 3.680 ;
        RECT  1.620 1.390 1.670 1.790 ;
        RECT  0.400 2.760 0.560 3.190 ;
        RECT  0.400 1.390 0.500 1.790 ;
        RECT  0.260 1.390 0.400 3.190 ;
        RECT  0.160 1.550 0.260 3.190 ;
    END
END INVX12

MACRO HOLDX1
    CLASS CORE ;
    FOREIGN HOLDX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION INOUT ;
        PORT
        LAYER met1 ;
        RECT  0.790 2.080 0.970 2.360 ;
        RECT  0.970 1.550 1.210 2.360 ;
        RECT  1.520 3.510 1.780 3.770 ;
        RECT  1.780 3.510 1.870 3.750 ;
        RECT  1.210 1.550 2.090 1.790 ;
        RECT  1.870 3.170 2.110 3.750 ;
        RECT  2.110 3.170 2.200 3.410 ;
        RECT  2.090 1.550 2.200 1.840 ;
        RECT  2.200 1.550 2.440 3.410 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 4.480 1.390 5.440 ;
        RECT  1.390 4.640 2.640 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.070 0.400 ;
        RECT  1.070 -0.400 1.080 0.930 ;
        RECT  1.080 -0.400 1.480 1.130 ;
        RECT  1.480 -0.400 1.490 0.930 ;
        RECT  1.490 -0.400 2.640 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.830 2.600 1.910 2.840 ;
        RECT  1.510 2.600 1.830 2.880 ;
        RECT  0.600 2.640 1.510 2.880 ;
        RECT  0.590 2.640 0.600 3.120 ;
        RECT  0.500 2.640 0.590 3.490 ;
        RECT  0.500 0.890 0.580 1.290 ;
        RECT  0.260 0.890 0.500 3.490 ;
        RECT  0.180 0.890 0.260 1.290 ;
        RECT  0.190 3.090 0.260 3.490 ;
    END
END HOLDX1

MACRO FILL8
    CLASS CORE ;
    FOREIGN FILL8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 5.280 0.400 ;
        END
    END GND
END FILL8

MACRO FILL64
    CLASS CORE ;
    FOREIGN FILL64 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 42.240 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 42.240 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 42.240 0.400 ;
        END
    END GND
END FILL64

MACRO FILL4
    CLASS CORE ;
    FOREIGN FILL4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 2.640 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 2.640 0.400 ;
        END
    END GND
END FILL4

MACRO FILL32
    CLASS CORE ;
    FOREIGN FILL32 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.120 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 21.120 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 21.120 0.400 ;
        END
    END GND
END FILL32

MACRO FILL2
    CLASS CORE ;
    FOREIGN FILL2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.320 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.320 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.320 0.400 ;
        END
    END GND
END FILL2

MACRO FILL16
    CLASS CORE ;
    FOREIGN FILL16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 10.560 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 10.560 0.400 ;
        END
    END GND
END FILL16

MACRO FILL1
    CLASS CORE ;
    FOREIGN FILL1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.660 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.660 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.660 0.400 ;
        END
    END GND
END FILL1

MACRO EDFFTRXL
    CLASS CORE ;
    FOREIGN EDFFTRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 3.940 2.150 4.370 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.230 3.620 16.710 3.860 ;
        RECT  16.700 2.390 16.710 2.650 ;
        RECT  16.480 1.320 16.710 2.070 ;
        RECT  16.710 1.320 16.720 3.860 ;
        RECT  16.720 1.830 16.950 3.860 ;
        RECT  16.950 2.390 16.960 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.710 3.480 14.720 4.320 ;
        RECT  14.720 3.480 14.870 4.330 ;
        RECT  14.870 3.100 14.980 4.330 ;
        RECT  14.980 3.100 15.110 4.320 ;
        RECT  15.160 0.720 15.560 1.100 ;
        RECT  15.110 3.100 15.960 3.340 ;
        RECT  15.560 0.860 15.960 1.100 ;
        RECT  15.960 0.860 16.200 3.340 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.820 1.860 2.840 2.100 ;
        RECT  2.840 1.830 3.100 2.100 ;
        RECT  3.100 1.860 5.160 2.100 ;
        RECT  5.160 1.860 5.560 2.200 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.880 2.380 6.060 2.620 ;
        RECT  6.060 1.840 6.140 2.620 ;
        RECT  6.140 1.830 6.300 2.620 ;
        RECT  6.300 1.830 6.400 2.090 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.700 2.000 0.770 2.400 ;
        RECT  0.770 0.720 0.860 2.400 ;
        RECT  0.860 0.710 1.010 2.400 ;
        RECT  1.010 0.710 1.120 0.970 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.760 5.440 ;
        RECT  0.760 4.480 1.160 5.440 ;
        RECT  1.160 4.640 4.180 5.440 ;
        RECT  4.180 4.480 4.620 5.440 ;
        RECT  4.620 4.640 8.060 5.440 ;
        RECT  8.060 4.480 8.460 5.440 ;
        RECT  8.460 4.640 10.540 5.440 ;
        RECT  10.540 4.480 10.940 5.440 ;
        RECT  10.940 4.640 13.280 5.440 ;
        RECT  13.280 3.210 13.520 5.440 ;
        RECT  13.520 4.640 15.470 5.440 ;
        RECT  15.470 3.650 15.870 5.440 ;
        RECT  15.870 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.540 0.400 ;
        RECT  1.540 -0.400 1.940 0.560 ;
        RECT  1.940 -0.400 8.370 0.400 ;
        RECT  8.370 -0.400 8.380 0.730 ;
        RECT  8.380 -0.400 8.780 0.850 ;
        RECT  8.780 -0.400 8.790 0.730 ;
        RECT  8.790 -0.400 11.750 0.400 ;
        RECT  11.750 -0.400 11.760 0.830 ;
        RECT  11.760 -0.400 12.160 0.950 ;
        RECT  12.160 -0.400 12.170 0.830 ;
        RECT  12.170 -0.400 14.390 0.400 ;
        RECT  14.390 -0.400 14.400 0.840 ;
        RECT  14.400 -0.400 14.800 1.040 ;
        RECT  14.800 -0.400 14.810 0.840 ;
        RECT  14.810 -0.400 16.490 0.400 ;
        RECT  16.490 -0.400 16.890 0.560 ;
        RECT  16.890 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  15.540 2.150 15.680 2.550 ;
        RECT  15.540 1.380 15.620 1.780 ;
        RECT  15.300 1.380 15.540 2.820 ;
        RECT  15.220 1.380 15.300 1.780 ;
        RECT  14.360 2.580 15.300 2.820 ;
        RECT  14.780 2.060 14.940 2.300 ;
        RECT  14.540 1.760 14.780 2.300 ;
        RECT  13.450 1.760 14.540 2.000 ;
        RECT  14.200 2.580 14.360 3.610 ;
        RECT  13.960 2.280 14.200 3.610 ;
        RECT  12.990 2.280 13.960 2.520 ;
        RECT  12.750 0.700 13.780 0.940 ;
        RECT  13.050 1.300 13.450 2.000 ;
        RECT  12.470 1.760 13.050 2.000 ;
        RECT  12.750 2.280 12.990 4.180 ;
        RECT  12.510 0.700 12.750 1.470 ;
        RECT  3.690 3.940 12.750 4.180 ;
        RECT  11.580 1.230 12.510 1.470 ;
        RECT  12.230 1.760 12.470 3.660 ;
        RECT  11.860 3.420 12.230 3.660 ;
        RECT  11.680 2.630 11.920 3.030 ;
        RECT  11.580 2.630 11.680 2.870 ;
        RECT  11.420 1.230 11.580 2.870 ;
        RECT  11.180 0.670 11.420 2.870 ;
        RECT  9.330 0.670 11.180 0.910 ;
        RECT  10.760 2.630 11.180 2.870 ;
        RECT  10.240 1.190 10.900 1.430 ;
        RECT  10.520 2.630 10.760 3.040 ;
        RECT  10.000 1.190 10.240 3.610 ;
        RECT  9.940 1.190 10.000 1.590 ;
        RECT  9.650 3.210 10.000 3.610 ;
        RECT  9.560 2.190 9.720 2.590 ;
        RECT  9.360 1.650 9.660 1.890 ;
        RECT  9.370 2.180 9.560 2.590 ;
        RECT  9.360 2.180 9.370 3.660 ;
        RECT  9.130 1.650 9.360 3.660 ;
        RECT  9.090 0.670 9.330 1.370 ;
        RECT  9.120 1.650 9.130 2.430 ;
        RECT  8.910 3.420 9.130 3.660 ;
        RECT  8.540 2.190 9.120 2.430 ;
        RECT  8.060 1.130 9.090 1.370 ;
        RECT  7.890 2.830 8.850 3.070 ;
        RECT  8.300 2.030 8.540 2.430 ;
        RECT  7.820 0.680 8.060 1.370 ;
        RECT  7.650 2.060 7.890 3.660 ;
        RECT  7.000 0.680 7.820 0.920 ;
        RECT  7.520 2.060 7.650 2.300 ;
        RECT  6.470 3.420 7.650 3.660 ;
        RECT  7.280 1.200 7.520 2.300 ;
        RECT  7.000 2.710 7.370 3.140 ;
        RECT  6.760 0.680 7.000 3.140 ;
        RECT  6.320 1.310 6.760 1.550 ;
        RECT  2.490 2.900 6.760 3.140 ;
        RECT  5.930 0.710 6.330 1.030 ;
        RECT  3.010 3.420 6.110 3.660 ;
        RECT  3.310 0.790 5.930 1.030 ;
        RECT  2.980 1.310 4.990 1.550 ;
        RECT  1.970 2.380 4.690 2.620 ;
        RECT  3.290 3.940 3.690 4.360 ;
        RECT  2.770 3.420 3.010 3.900 ;
        RECT  2.740 0.640 2.980 1.550 ;
        RECT  2.570 0.640 2.740 0.880 ;
        RECT  2.250 2.900 2.490 3.670 ;
        RECT  0.570 3.430 2.250 3.670 ;
        RECT  1.540 1.290 2.110 1.530 ;
        RECT  1.730 2.380 1.970 3.150 ;
        RECT  1.540 2.380 1.730 2.620 ;
        RECT  1.300 1.290 1.540 2.620 ;
        RECT  0.420 2.750 0.570 3.670 ;
        RECT  0.420 1.170 0.490 1.610 ;
        RECT  0.330 1.170 0.420 3.670 ;
        RECT  0.180 1.170 0.330 3.150 ;
        RECT  0.170 2.750 0.180 3.150 ;
    END
END EDFFTRXL

MACRO EDFFTRX4
    CLASS CORE ;
    FOREIGN EDFFTRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ EDFFTRXL ;
    SIZE 21.780 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.510 3.780 1.930 4.340 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  19.910 1.260 19.930 2.660 ;
        RECT  19.930 1.260 20.350 3.180 ;
        RECT  20.350 2.760 20.520 3.180 ;
        RECT  20.350 1.270 20.600 1.670 ;
        RECT  20.520 2.770 20.720 3.170 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.590 1.260 18.610 2.660 ;
        RECT  18.610 1.260 19.030 3.180 ;
        RECT  19.030 1.260 19.040 2.170 ;
        RECT  19.030 2.770 19.180 3.170 ;
        RECT  19.040 1.270 19.180 1.670 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.030 1.850 2.840 2.090 ;
        RECT  2.840 1.830 2.970 2.090 ;
        RECT  2.970 1.820 5.080 2.100 ;
        RECT  5.080 1.750 5.370 2.100 ;
        RECT  5.370 1.740 5.650 2.100 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.320 4.020 6.140 4.260 ;
        RECT  6.140 4.020 6.390 4.330 ;
        RECT  6.390 4.070 6.400 4.330 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 1.950 0.780 2.350 ;
        RECT  0.780 1.840 0.860 2.350 ;
        RECT  0.860 1.830 1.020 2.350 ;
        RECT  1.020 1.830 1.120 2.090 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.860 5.440 ;
        RECT  0.860 3.940 1.100 5.440 ;
        RECT  1.100 4.640 2.210 5.440 ;
        RECT  2.210 3.910 2.220 5.440 ;
        RECT  2.220 3.790 2.620 5.440 ;
        RECT  2.620 3.910 2.630 5.440 ;
        RECT  2.630 4.640 4.280 5.440 ;
        RECT  4.280 4.050 4.290 5.440 ;
        RECT  4.290 3.930 4.690 5.440 ;
        RECT  4.690 4.050 4.700 5.440 ;
        RECT  4.700 4.640 7.880 5.440 ;
        RECT  7.880 4.480 8.860 5.440 ;
        RECT  8.860 4.640 11.330 5.440 ;
        RECT  11.330 4.480 11.730 5.440 ;
        RECT  11.730 4.640 13.890 5.440 ;
        RECT  13.890 4.480 14.290 5.440 ;
        RECT  14.290 4.640 16.500 5.440 ;
        RECT  16.500 4.480 16.900 5.440 ;
        RECT  16.900 4.640 18.040 5.440 ;
        RECT  18.040 4.030 18.440 5.440 ;
        RECT  18.440 4.640 19.590 5.440 ;
        RECT  19.590 4.230 19.600 5.440 ;
        RECT  19.600 4.030 20.000 5.440 ;
        RECT  20.000 4.230 20.010 5.440 ;
        RECT  20.010 4.640 20.980 5.440 ;
        RECT  20.980 4.230 20.990 5.440 ;
        RECT  20.990 4.030 21.390 5.440 ;
        RECT  21.390 4.230 21.400 5.440 ;
        RECT  21.400 4.640 21.780 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 2.090 0.400 ;
        RECT  2.090 -0.400 2.490 0.560 ;
        RECT  2.490 -0.400 8.650 0.400 ;
        RECT  8.650 -0.400 8.660 1.110 ;
        RECT  8.660 -0.400 9.060 1.230 ;
        RECT  9.060 -0.400 9.070 1.110 ;
        RECT  9.070 -0.400 10.170 0.400 ;
        RECT  10.170 -0.400 10.180 1.110 ;
        RECT  10.180 -0.400 10.580 1.230 ;
        RECT  10.580 -0.400 10.590 1.110 ;
        RECT  10.590 -0.400 11.880 0.400 ;
        RECT  11.880 -0.400 11.890 0.930 ;
        RECT  11.890 -0.400 12.290 1.130 ;
        RECT  12.290 -0.400 12.300 0.930 ;
        RECT  12.300 -0.400 14.320 0.400 ;
        RECT  14.320 -0.400 14.330 0.720 ;
        RECT  14.330 -0.400 14.730 0.840 ;
        RECT  14.730 -0.400 14.740 0.720 ;
        RECT  14.740 -0.400 16.770 0.400 ;
        RECT  16.770 -0.400 17.170 0.560 ;
        RECT  17.170 -0.400 18.100 0.400 ;
        RECT  18.100 -0.400 18.110 0.790 ;
        RECT  18.110 -0.400 18.510 0.990 ;
        RECT  18.510 -0.400 18.520 0.790 ;
        RECT  18.520 -0.400 19.530 0.400 ;
        RECT  19.530 -0.400 19.540 0.790 ;
        RECT  19.540 -0.400 19.940 0.990 ;
        RECT  19.940 -0.400 19.950 0.790 ;
        RECT  19.950 -0.400 20.860 0.400 ;
        RECT  20.860 -0.400 20.870 0.790 ;
        RECT  20.870 -0.400 21.270 0.990 ;
        RECT  21.270 -0.400 21.280 0.790 ;
        RECT  21.280 -0.400 21.780 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  21.020 2.200 21.260 3.720 ;
        RECT  18.320 3.480 21.020 3.720 ;
        RECT  18.080 1.430 18.320 3.720 ;
        RECT  17.900 1.430 18.080 1.670 ;
        RECT  17.560 2.910 18.080 3.310 ;
        RECT  17.500 1.270 17.900 1.670 ;
        RECT  17.610 1.970 17.800 2.370 ;
        RECT  17.040 1.970 17.610 2.380 ;
        RECT  17.320 2.910 17.560 4.180 ;
        RECT  16.340 3.940 17.320 4.180 ;
        RECT  16.800 1.170 17.040 3.660 ;
        RECT  15.950 1.170 16.800 1.410 ;
        RECT  12.610 3.420 16.800 3.660 ;
        RECT  16.330 1.990 16.490 2.390 ;
        RECT  15.940 3.940 16.340 4.240 ;
        RECT  16.090 1.990 16.330 3.140 ;
        RECT  15.330 2.900 16.090 3.140 ;
        RECT  15.630 1.120 15.950 1.410 ;
        RECT  7.310 3.940 15.940 4.180 ;
        RECT  15.370 1.690 15.770 2.090 ;
        RECT  13.510 1.120 15.630 1.360 ;
        RECT  14.440 1.690 15.370 1.930 ;
        RECT  14.860 2.680 15.330 3.140 ;
        RECT  13.250 2.900 14.860 3.140 ;
        RECT  13.990 2.370 14.620 2.610 ;
        RECT  14.200 1.640 14.440 1.930 ;
        RECT  12.800 1.640 14.200 1.880 ;
        RECT  13.720 2.160 13.990 2.610 ;
        RECT  12.340 2.160 13.720 2.400 ;
        RECT  13.110 0.740 13.510 1.360 ;
        RECT  12.850 2.680 13.250 3.140 ;
        RECT  11.510 2.900 12.850 3.140 ;
        RECT  12.560 1.560 12.800 1.880 ;
        RECT  11.530 1.560 12.560 1.800 ;
        RECT  12.310 2.080 12.340 2.400 ;
        RECT  11.910 2.080 12.310 2.480 ;
        RECT  10.990 2.080 11.910 2.320 ;
        RECT  11.130 0.880 11.530 1.800 ;
        RECT  11.270 2.600 11.510 3.660 ;
        RECT  9.130 3.420 11.270 3.660 ;
        RECT  10.470 1.560 11.130 1.800 ;
        RECT  10.750 2.080 10.990 3.140 ;
        RECT  9.650 2.900 10.750 3.140 ;
        RECT  10.230 1.560 10.470 2.620 ;
        RECT  10.070 2.380 10.230 2.620 ;
        RECT  9.650 0.990 9.820 1.230 ;
        RECT  9.410 0.990 9.650 3.140 ;
        RECT  8.720 1.510 9.410 1.770 ;
        RECT  8.890 2.190 9.130 3.660 ;
        RECT  8.200 2.190 8.890 2.430 ;
        RECT  8.480 1.510 8.720 1.910 ;
        RECT  7.680 2.720 8.610 2.960 ;
        RECT  7.960 0.670 8.200 2.430 ;
        RECT  7.050 0.670 7.960 0.910 ;
        RECT  7.570 1.350 7.680 3.660 ;
        RECT  7.440 1.190 7.570 3.660 ;
        RECT  7.330 1.190 7.440 1.590 ;
        RECT  6.520 3.420 7.440 3.660 ;
        RECT  6.910 3.940 7.310 4.370 ;
        RECT  7.050 2.540 7.160 2.940 ;
        RECT  6.810 0.670 7.050 3.130 ;
        RECT  6.450 1.400 6.810 1.640 ;
        RECT  2.540 2.890 6.810 3.130 ;
        RECT  6.290 0.670 6.530 1.120 ;
        RECT  3.650 0.670 6.290 0.910 ;
        RECT  3.400 3.410 5.970 3.650 ;
        RECT  3.310 1.190 5.330 1.430 ;
        RECT  2.020 2.370 4.830 2.610 ;
        RECT  3.000 3.410 3.400 3.860 ;
        RECT  3.070 0.720 3.310 1.430 ;
        RECT  2.910 0.720 3.070 1.120 ;
        RECT  2.300 2.890 2.540 3.510 ;
        RECT  0.570 3.270 2.300 3.510 ;
        RECT  1.860 2.370 2.020 2.990 ;
        RECT  1.750 2.360 1.860 2.990 ;
        RECT  1.510 1.230 1.750 2.990 ;
        RECT  0.400 2.750 0.570 3.510 ;
        RECT  0.400 1.310 0.490 1.710 ;
        RECT  0.330 1.310 0.400 3.510 ;
        RECT  0.160 1.310 0.330 3.150 ;
    END
END EDFFTRX4

MACRO EDFFTRX2
    CLASS CORE ;
    FOREIGN EDFFTRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ EDFFTRXL ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 4.070 1.780 4.330 ;
        RECT  1.780 4.080 2.490 4.320 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.360 3.510 17.470 3.770 ;
        RECT  17.470 3.500 17.620 3.770 ;
        RECT  17.620 3.500 17.920 3.780 ;
        RECT  17.420 0.760 17.920 1.000 ;
        RECT  17.920 0.760 18.040 3.780 ;
        RECT  18.040 0.760 18.160 3.740 ;
        RECT  18.160 3.060 18.320 3.520 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.780 0.720 16.180 1.120 ;
        RECT  16.180 0.880 16.400 1.120 ;
        RECT  16.400 0.880 16.640 1.520 ;
        RECT  16.440 2.950 16.810 3.950 ;
        RECT  16.810 2.490 16.840 3.950 ;
        RECT  16.840 2.490 16.960 3.210 ;
        RECT  16.960 2.490 17.050 3.190 ;
        RECT  17.050 2.490 17.420 2.730 ;
        RECT  16.640 1.280 17.420 1.520 ;
        RECT  17.420 1.280 17.660 2.730 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.820 1.860 2.840 2.100 ;
        RECT  2.840 1.830 3.100 2.100 ;
        RECT  3.100 1.860 5.560 2.100 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.840 2.220 6.000 2.620 ;
        RECT  6.000 1.850 6.140 2.620 ;
        RECT  6.140 1.830 6.240 2.620 ;
        RECT  6.240 1.830 6.400 2.090 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.000 0.770 2.400 ;
        RECT  0.770 0.720 0.860 2.400 ;
        RECT  0.860 0.710 1.010 2.400 ;
        RECT  1.010 0.710 1.120 0.970 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.760 5.440 ;
        RECT  0.760 4.480 1.160 5.440 ;
        RECT  1.160 4.640 4.180 5.440 ;
        RECT  4.180 4.480 4.620 5.440 ;
        RECT  4.620 4.640 8.060 5.440 ;
        RECT  8.060 4.480 8.460 5.440 ;
        RECT  8.460 4.640 10.560 5.440 ;
        RECT  10.560 4.480 10.960 5.440 ;
        RECT  10.960 4.640 13.140 5.440 ;
        RECT  13.140 4.480 13.540 5.440 ;
        RECT  13.540 4.640 14.930 5.440 ;
        RECT  14.930 3.480 14.940 5.440 ;
        RECT  14.940 3.280 15.340 5.440 ;
        RECT  15.340 3.480 15.350 5.440 ;
        RECT  15.350 4.640 17.260 5.440 ;
        RECT  17.260 4.150 17.660 5.440 ;
        RECT  17.660 4.640 18.480 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.480 0.400 ;
        RECT  1.480 -0.400 1.880 0.560 ;
        RECT  1.880 -0.400 8.370 0.400 ;
        RECT  8.370 -0.400 8.380 0.730 ;
        RECT  8.380 -0.400 8.780 0.850 ;
        RECT  8.780 -0.400 8.790 0.730 ;
        RECT  8.790 -0.400 11.760 0.400 ;
        RECT  11.760 -0.400 12.180 1.320 ;
        RECT  12.180 -0.400 14.430 0.400 ;
        RECT  14.430 -0.400 14.830 0.560 ;
        RECT  14.830 -0.400 16.600 0.400 ;
        RECT  16.600 -0.400 17.000 0.560 ;
        RECT  17.000 -0.400 18.480 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.100 1.800 17.130 2.200 ;
        RECT  15.860 1.400 16.100 3.520 ;
        RECT  15.440 1.400 15.860 1.640 ;
        RECT  15.700 2.760 15.860 3.520 ;
        RECT  14.630 2.760 15.700 3.000 ;
        RECT  15.340 1.920 15.580 2.480 ;
        RECT  15.040 1.190 15.440 1.640 ;
        RECT  13.490 1.920 15.340 2.160 ;
        RECT  14.390 2.760 14.630 4.310 ;
        RECT  14.230 3.940 14.390 4.310 ;
        RECT  12.840 3.940 14.230 4.180 ;
        RECT  13.330 3.210 14.000 3.660 ;
        RECT  12.810 0.700 13.820 0.940 ;
        RECT  13.330 1.430 13.490 2.160 ;
        RECT  13.090 1.430 13.330 3.660 ;
        RECT  12.260 3.420 13.090 3.660 ;
        RECT  12.600 3.940 12.840 4.360 ;
        RECT  12.570 0.700 12.810 2.030 ;
        RECT  11.580 4.120 12.600 4.360 ;
        RECT  11.480 1.790 12.570 2.030 ;
        RECT  11.860 3.420 12.260 3.830 ;
        RECT  11.620 2.730 12.020 3.140 ;
        RECT  11.480 2.730 11.620 2.970 ;
        RECT  11.340 3.940 11.580 4.360 ;
        RECT  11.420 1.790 11.480 2.970 ;
        RECT  11.180 0.670 11.420 2.970 ;
        RECT  3.690 3.940 11.340 4.180 ;
        RECT  9.330 0.670 11.180 0.910 ;
        RECT  10.760 2.730 11.180 2.970 ;
        RECT  10.240 1.190 10.900 1.430 ;
        RECT  10.520 2.730 10.760 3.140 ;
        RECT  10.000 1.190 10.240 3.660 ;
        RECT  9.650 3.420 10.000 3.660 ;
        RECT  9.480 1.650 9.720 3.140 ;
        RECT  9.260 1.650 9.480 2.180 ;
        RECT  9.370 2.900 9.480 3.140 ;
        RECT  9.130 2.900 9.370 3.570 ;
        RECT  9.090 0.670 9.330 1.370 ;
        RECT  8.540 1.940 9.260 2.180 ;
        RECT  8.730 3.330 9.130 3.570 ;
        RECT  8.060 1.130 9.090 1.370 ;
        RECT  7.890 2.750 8.830 2.990 ;
        RECT  8.300 1.940 8.540 2.340 ;
        RECT  7.820 0.680 8.060 1.370 ;
        RECT  7.650 2.060 7.890 3.660 ;
        RECT  7.000 0.680 7.820 0.920 ;
        RECT  7.520 2.060 7.650 2.300 ;
        RECT  6.470 3.420 7.650 3.660 ;
        RECT  7.280 1.200 7.520 2.300 ;
        RECT  7.000 2.710 7.370 3.140 ;
        RECT  6.760 0.680 7.000 3.140 ;
        RECT  6.470 1.310 6.760 1.550 ;
        RECT  2.490 2.900 6.760 3.140 ;
        RECT  6.030 0.730 6.430 1.030 ;
        RECT  3.010 3.420 6.050 3.660 ;
        RECT  3.250 0.790 6.030 1.030 ;
        RECT  2.910 1.310 4.990 1.550 ;
        RECT  1.970 2.380 4.580 2.620 ;
        RECT  3.290 3.940 3.690 4.270 ;
        RECT  2.770 3.420 3.010 3.830 ;
        RECT  2.670 0.670 2.910 1.550 ;
        RECT  2.510 0.670 2.670 0.910 ;
        RECT  2.250 2.900 2.490 3.670 ;
        RECT  0.490 3.430 2.250 3.670 ;
        RECT  1.540 1.250 2.050 1.490 ;
        RECT  1.730 2.380 1.970 3.150 ;
        RECT  1.540 2.380 1.730 2.620 ;
        RECT  1.300 1.250 1.540 2.620 ;
        RECT  0.400 1.170 0.490 1.570 ;
        RECT  0.400 2.920 0.490 3.670 ;
        RECT  0.250 1.170 0.400 3.670 ;
        RECT  0.160 1.170 0.250 3.240 ;
    END
END EDFFTRX2

MACRO EDFFTRX1
    CLASS CORE ;
    FOREIGN EDFFTRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ EDFFTRXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 4.070 1.530 4.330 ;
        RECT  1.530 4.010 1.780 4.330 ;
        RECT  1.780 4.010 2.490 4.250 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.230 3.620 16.520 4.020 ;
        RECT  16.520 3.620 16.710 4.030 ;
        RECT  16.700 2.390 16.710 2.650 ;
        RECT  16.480 1.320 16.710 2.070 ;
        RECT  16.710 1.320 16.720 4.030 ;
        RECT  16.720 1.830 16.950 4.030 ;
        RECT  16.950 3.650 16.960 4.030 ;
        RECT  16.950 2.390 16.960 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.710 3.480 14.870 3.880 ;
        RECT  14.870 3.100 15.110 3.880 ;
        RECT  15.160 0.670 15.560 1.100 ;
        RECT  15.110 3.100 15.960 3.340 ;
        RECT  15.560 0.860 15.960 1.100 ;
        RECT  15.960 0.860 16.200 3.340 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.820 1.860 2.840 2.100 ;
        RECT  2.840 1.830 3.100 2.100 ;
        RECT  3.100 1.860 4.910 2.100 ;
        RECT  4.910 1.860 5.310 2.120 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.480 1.270 5.590 1.530 ;
        RECT  5.590 1.270 5.740 2.350 ;
        RECT  5.740 1.280 5.830 2.350 ;
        RECT  5.830 1.950 5.950 2.350 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.000 0.770 2.400 ;
        RECT  0.770 0.720 0.860 2.400 ;
        RECT  0.860 0.710 0.920 2.400 ;
        RECT  0.920 0.710 1.010 2.320 ;
        RECT  1.010 0.710 1.120 0.970 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.760 5.440 ;
        RECT  0.760 4.480 1.160 5.440 ;
        RECT  1.160 4.640 4.110 5.440 ;
        RECT  4.110 4.480 4.510 5.440 ;
        RECT  4.510 4.640 7.820 5.440 ;
        RECT  7.820 4.480 8.220 5.440 ;
        RECT  8.220 4.640 10.530 5.440 ;
        RECT  10.530 4.480 10.930 5.440 ;
        RECT  10.930 4.640 13.280 5.440 ;
        RECT  13.280 3.280 13.520 5.440 ;
        RECT  13.520 4.640 15.470 5.440 ;
        RECT  15.470 3.700 15.870 5.440 ;
        RECT  15.870 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.480 0.400 ;
        RECT  1.480 -0.400 1.880 0.560 ;
        RECT  1.880 -0.400 8.370 0.400 ;
        RECT  8.370 -0.400 8.380 0.730 ;
        RECT  8.380 -0.400 8.780 0.850 ;
        RECT  8.780 -0.400 8.790 0.730 ;
        RECT  8.790 -0.400 11.760 0.400 ;
        RECT  11.760 -0.400 11.770 0.830 ;
        RECT  11.770 -0.400 12.170 0.950 ;
        RECT  12.170 -0.400 12.180 0.830 ;
        RECT  12.180 -0.400 14.390 0.400 ;
        RECT  14.390 -0.400 14.400 0.760 ;
        RECT  14.400 -0.400 14.800 0.960 ;
        RECT  14.800 -0.400 14.810 0.760 ;
        RECT  14.810 -0.400 16.480 0.400 ;
        RECT  16.480 -0.400 16.880 0.560 ;
        RECT  16.880 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  15.620 2.150 15.680 2.550 ;
        RECT  15.300 1.380 15.620 2.820 ;
        RECT  15.220 1.380 15.300 1.780 ;
        RECT  14.260 2.580 15.300 2.820 ;
        RECT  14.780 2.060 14.940 2.300 ;
        RECT  14.540 1.760 14.780 2.300 ;
        RECT  13.450 1.760 14.540 2.000 ;
        RECT  14.260 3.290 14.360 3.690 ;
        RECT  14.020 2.280 14.260 3.690 ;
        RECT  12.990 2.280 14.020 2.520 ;
        RECT  13.960 3.290 14.020 3.690 ;
        RECT  12.750 0.700 13.780 0.940 ;
        RECT  13.050 1.300 13.450 2.000 ;
        RECT  12.470 1.760 13.050 2.000 ;
        RECT  12.750 2.280 12.990 4.180 ;
        RECT  12.510 0.700 12.750 1.470 ;
        RECT  3.290 3.940 12.750 4.180 ;
        RECT  11.580 1.230 12.510 1.470 ;
        RECT  12.230 1.760 12.470 3.660 ;
        RECT  11.860 3.420 12.230 3.660 ;
        RECT  11.680 2.630 11.920 3.030 ;
        RECT  11.580 2.630 11.680 2.870 ;
        RECT  11.420 1.230 11.580 2.870 ;
        RECT  11.260 0.670 11.420 2.870 ;
        RECT  11.180 0.670 11.260 1.870 ;
        RECT  10.760 2.630 11.260 2.870 ;
        RECT  9.330 0.670 11.180 0.910 ;
        RECT  10.240 1.190 10.900 1.430 ;
        RECT  10.520 2.630 10.760 3.040 ;
        RECT  10.000 1.190 10.240 3.530 ;
        RECT  9.940 1.190 10.000 1.590 ;
        RECT  9.650 3.290 10.000 3.530 ;
        RECT  9.660 2.190 9.720 2.590 ;
        RECT  9.370 1.650 9.660 2.590 ;
        RECT  9.260 1.650 9.370 3.660 ;
        RECT  9.090 0.670 9.330 1.370 ;
        RECT  9.130 2.190 9.260 3.660 ;
        RECT  8.490 2.190 9.130 2.430 ;
        RECT  8.730 3.420 9.130 3.660 ;
        RECT  7.890 1.130 9.090 1.370 ;
        RECT  7.630 2.830 8.830 3.070 ;
        RECT  8.090 2.030 8.490 2.430 ;
        RECT  7.650 0.680 7.890 1.370 ;
        RECT  6.850 0.680 7.650 0.920 ;
        RECT  7.390 2.060 7.630 3.660 ;
        RECT  7.370 2.060 7.390 2.300 ;
        RECT  6.470 3.420 7.390 3.660 ;
        RECT  7.130 1.200 7.370 2.300 ;
        RECT  6.850 2.710 7.110 3.140 ;
        RECT  6.610 0.680 6.850 3.140 ;
        RECT  6.320 1.310 6.610 1.550 ;
        RECT  2.490 2.900 6.610 3.140 ;
        RECT  3.650 0.720 6.330 0.960 ;
        RECT  3.010 3.420 5.990 3.660 ;
        RECT  2.910 1.310 4.990 1.550 ;
        RECT  1.970 2.380 4.580 2.620 ;
        RECT  3.250 0.720 3.650 1.030 ;
        RECT  2.770 3.420 3.010 3.820 ;
        RECT  2.670 0.670 2.910 1.550 ;
        RECT  2.510 0.670 2.670 0.910 ;
        RECT  2.250 2.900 2.490 3.670 ;
        RECT  0.570 3.430 2.250 3.670 ;
        RECT  1.540 1.250 2.050 1.490 ;
        RECT  1.730 2.380 1.970 3.150 ;
        RECT  1.540 2.380 1.730 2.620 ;
        RECT  1.300 1.250 1.540 2.620 ;
        RECT  0.400 2.760 0.570 3.670 ;
        RECT  0.400 1.170 0.490 1.570 ;
        RECT  0.330 1.170 0.400 3.670 ;
        RECT  0.170 1.170 0.330 3.160 ;
        RECT  0.160 1.170 0.170 3.080 ;
    END
END EDFFTRX1

MACRO EDFFXL
    CLASS CORE ;
    FOREIGN EDFFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.610 2.840 14.630 3.240 ;
        RECT  14.610 1.400 14.720 1.960 ;
        RECT  14.630 2.520 14.730 3.240 ;
        RECT  14.720 1.400 14.730 2.090 ;
        RECT  14.730 1.400 14.970 3.240 ;
        RECT  14.970 1.400 14.980 2.090 ;
        RECT  14.970 2.520 15.010 3.240 ;
        RECT  14.980 1.400 15.010 1.960 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.990 3.630 13.150 4.030 ;
        RECT  13.150 3.530 13.390 4.030 ;
        RECT  12.990 0.730 13.390 1.100 ;
        RECT  13.390 3.530 13.400 3.770 ;
        RECT  13.400 3.510 13.660 3.770 ;
        RECT  13.660 3.510 14.090 3.750 ;
        RECT  13.390 0.860 14.090 1.100 ;
        RECT  14.090 0.860 14.330 3.750 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 3.960 2.000 4.360 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.530 2.130 4.730 2.370 ;
        RECT  4.730 2.130 4.820 2.630 ;
        RECT  4.820 2.130 4.970 2.650 ;
        RECT  4.970 2.390 5.080 2.650 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.690 2.090 0.860 2.640 ;
        RECT  0.860 2.090 0.930 2.650 ;
        RECT  0.930 2.390 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.780 5.440 ;
        RECT  0.780 4.480 1.180 5.440 ;
        RECT  1.180 4.640 3.730 5.440 ;
        RECT  3.730 4.480 4.130 5.440 ;
        RECT  4.130 4.640 7.280 5.440 ;
        RECT  7.280 4.480 7.680 5.440 ;
        RECT  7.680 4.640 8.880 5.440 ;
        RECT  8.880 4.480 9.860 5.440 ;
        RECT  9.860 4.640 12.170 5.440 ;
        RECT  12.170 4.480 12.570 5.440 ;
        RECT  12.570 4.640 13.790 5.440 ;
        RECT  13.790 4.480 14.190 5.440 ;
        RECT  14.190 4.640 15.180 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.950 0.400 ;
        RECT  0.950 -0.400 1.350 0.560 ;
        RECT  1.350 -0.400 3.400 0.400 ;
        RECT  3.400 -0.400 3.800 0.560 ;
        RECT  3.800 -0.400 6.950 0.400 ;
        RECT  6.950 -0.400 6.960 1.070 ;
        RECT  6.960 -0.400 7.360 1.270 ;
        RECT  7.360 -0.400 7.370 1.070 ;
        RECT  7.370 -0.400 9.570 0.400 ;
        RECT  9.570 -0.400 9.580 0.800 ;
        RECT  9.580 -0.400 9.980 1.000 ;
        RECT  9.980 -0.400 9.990 0.800 ;
        RECT  9.990 -0.400 12.110 0.400 ;
        RECT  12.110 -0.400 12.510 0.560 ;
        RECT  12.510 -0.400 13.730 0.400 ;
        RECT  13.730 -0.400 14.130 0.560 ;
        RECT  14.130 -0.400 15.180 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  13.570 1.550 13.810 3.010 ;
        RECT  13.390 1.550 13.570 1.790 ;
        RECT  13.450 2.770 13.570 3.010 ;
        RECT  13.050 2.770 13.450 3.170 ;
        RECT  12.990 1.390 13.390 1.790 ;
        RECT  11.890 2.930 13.050 3.170 ;
        RECT  12.470 2.070 12.870 2.470 ;
        RECT  11.310 2.150 12.470 2.390 ;
        RECT  11.650 2.930 11.890 4.340 ;
        RECT  11.490 3.940 11.650 4.340 ;
        RECT  10.590 0.760 11.590 1.000 ;
        RECT  3.090 3.940 11.490 4.180 ;
        RECT  11.180 1.440 11.310 3.660 ;
        RECT  11.070 1.280 11.180 3.660 ;
        RECT  10.940 1.280 11.070 1.680 ;
        RECT  10.890 3.260 11.070 3.660 ;
        RECT  10.590 2.580 10.790 2.980 ;
        RECT  10.350 0.760 10.590 3.660 ;
        RECT  5.950 3.420 10.350 3.660 ;
        RECT  9.830 1.560 10.070 3.140 ;
        RECT  9.160 1.560 9.830 1.800 ;
        RECT  8.990 2.900 9.830 3.140 ;
        RECT  8.550 2.330 9.550 2.570 ;
        RECT  8.920 0.670 9.160 1.800 ;
        RECT  8.680 0.670 8.920 0.910 ;
        RECT  8.470 2.330 8.550 3.060 ;
        RECT  8.240 1.550 8.470 3.060 ;
        RECT  8.230 0.910 8.240 3.060 ;
        RECT  7.840 0.910 8.230 1.790 ;
        RECT  8.150 2.820 8.230 3.060 ;
        RECT  7.710 2.140 7.950 2.540 ;
        RECT  6.990 1.550 7.840 1.790 ;
        RECT  6.470 2.300 7.710 2.540 ;
        RECT  6.750 1.550 6.990 2.020 ;
        RECT  6.230 1.080 6.470 3.140 ;
        RECT  6.020 1.080 6.230 1.320 ;
        RECT  5.620 0.920 6.020 1.320 ;
        RECT  5.710 1.600 5.950 3.660 ;
        RECT  2.740 1.600 5.710 1.840 ;
        RECT  5.190 3.200 5.430 3.660 ;
        RECT  2.450 3.420 5.190 3.660 ;
        RECT  4.980 0.920 5.140 1.320 ;
        RECT  4.740 0.860 4.980 1.320 ;
        RECT  2.460 0.860 4.740 1.100 ;
        RECT  3.300 2.850 4.460 3.090 ;
        RECT  3.060 2.140 3.300 3.090 ;
        RECT  2.690 3.940 3.090 4.270 ;
        RECT  2.110 2.140 3.060 2.380 ;
        RECT  2.500 1.380 2.740 1.840 ;
        RECT  0.570 1.380 2.500 1.620 ;
        RECT  2.060 0.790 2.460 1.100 ;
        RECT  2.050 1.900 2.110 2.380 ;
        RECT  1.810 1.900 2.050 3.680 ;
        RECT  1.710 1.900 1.810 2.140 ;
        RECT  1.650 3.280 1.810 3.680 ;
        RECT  0.410 1.290 0.570 1.690 ;
        RECT  0.410 3.280 0.570 3.680 ;
        RECT  0.170 1.290 0.410 3.680 ;
    END
END EDFFXL

MACRO EDFFX4
    CLASS CORE ;
    FOREIGN EDFFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ EDFFXL ;
    SIZE 20.460 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  19.220 2.870 19.250 3.270 ;
        RECT  19.220 1.250 19.250 1.650 ;
        RECT  19.250 1.250 19.620 3.270 ;
        RECT  19.620 1.260 19.650 3.270 ;
        RECT  19.650 1.260 19.690 2.660 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.680 2.870 17.930 3.270 ;
        RECT  17.880 1.250 17.930 1.650 ;
        RECT  17.930 1.250 18.280 3.270 ;
        RECT  18.280 1.260 18.330 3.270 ;
        RECT  18.330 1.260 18.370 2.660 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.420 1.590 3.430 2.090 ;
        RECT  3.430 1.470 3.830 2.090 ;
        RECT  3.830 1.590 3.840 2.090 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.480 1.460 4.730 1.860 ;
        RECT  4.730 1.460 4.820 2.080 ;
        RECT  4.820 1.460 4.880 2.090 ;
        RECT  4.880 1.620 4.970 2.090 ;
        RECT  4.970 1.830 5.080 2.090 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.360 2.650 ;
        RECT  0.360 2.060 0.460 2.650 ;
        RECT  0.460 2.060 0.600 2.630 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.040 5.440 ;
        RECT  1.040 4.480 1.440 5.440 ;
        RECT  1.440 4.640 3.600 5.440 ;
        RECT  3.600 4.480 4.000 5.440 ;
        RECT  4.000 4.640 7.260 5.440 ;
        RECT  7.260 4.480 7.660 5.440 ;
        RECT  7.660 4.640 9.780 5.440 ;
        RECT  9.780 4.480 10.180 5.440 ;
        RECT  10.180 4.640 12.630 5.440 ;
        RECT  12.630 4.480 13.030 5.440 ;
        RECT  13.030 4.640 15.430 5.440 ;
        RECT  15.430 4.480 15.830 5.440 ;
        RECT  15.830 4.640 16.970 5.440 ;
        RECT  16.970 4.320 16.980 5.440 ;
        RECT  16.980 4.120 17.380 5.440 ;
        RECT  17.380 4.320 17.390 5.440 ;
        RECT  17.390 4.640 18.480 5.440 ;
        RECT  18.480 4.330 18.490 5.440 ;
        RECT  18.490 4.130 18.890 5.440 ;
        RECT  18.890 4.330 18.900 5.440 ;
        RECT  18.900 4.640 19.880 5.440 ;
        RECT  19.880 4.350 19.890 5.440 ;
        RECT  19.890 4.150 20.290 5.440 ;
        RECT  20.290 4.350 20.300 5.440 ;
        RECT  20.300 4.640 20.460 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.920 0.400 ;
        RECT  0.920 -0.400 0.930 0.730 ;
        RECT  0.930 -0.400 1.330 0.930 ;
        RECT  1.330 -0.400 1.340 0.730 ;
        RECT  1.340 -0.400 3.180 0.400 ;
        RECT  3.180 -0.400 3.640 0.560 ;
        RECT  3.640 -0.400 6.830 0.400 ;
        RECT  6.830 -0.400 6.840 1.010 ;
        RECT  6.840 -0.400 7.240 1.130 ;
        RECT  7.240 -0.400 7.250 1.010 ;
        RECT  7.250 -0.400 8.620 0.400 ;
        RECT  8.620 -0.400 8.860 1.330 ;
        RECT  8.860 -0.400 10.490 0.400 ;
        RECT  10.490 -0.400 10.890 0.560 ;
        RECT  10.890 -0.400 13.050 0.400 ;
        RECT  13.050 -0.400 13.450 0.560 ;
        RECT  13.450 -0.400 15.830 0.400 ;
        RECT  15.830 -0.400 16.230 1.610 ;
        RECT  16.230 -0.400 17.270 0.400 ;
        RECT  17.270 -0.400 17.670 0.970 ;
        RECT  17.670 -0.400 18.540 0.400 ;
        RECT  18.540 -0.400 18.550 0.770 ;
        RECT  18.550 -0.400 18.950 0.970 ;
        RECT  18.950 -0.400 18.960 0.770 ;
        RECT  18.960 -0.400 19.880 0.400 ;
        RECT  19.880 -0.400 19.890 0.770 ;
        RECT  19.890 -0.400 20.290 0.970 ;
        RECT  20.290 -0.400 20.300 0.770 ;
        RECT  20.300 -0.400 20.460 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  19.930 2.260 20.170 3.840 ;
        RECT  17.440 3.600 19.930 3.840 ;
        RECT  17.200 1.220 17.440 3.840 ;
        RECT  16.950 1.220 17.200 1.460 ;
        RECT  16.170 3.440 17.200 3.840 ;
        RECT  15.580 1.940 16.960 2.340 ;
        RECT  16.550 1.060 16.950 1.460 ;
        RECT  15.930 2.660 16.170 4.180 ;
        RECT  12.010 3.940 15.930 4.180 ;
        RECT  15.340 1.260 15.580 3.660 ;
        RECT  15.020 1.260 15.340 1.500 ;
        RECT  11.670 3.420 15.340 3.660 ;
        RECT  14.860 1.860 15.100 2.850 ;
        RECT  14.780 0.950 15.020 1.500 ;
        RECT  14.050 2.610 14.860 2.850 ;
        RECT  14.740 0.950 14.780 1.190 ;
        RECT  14.340 0.790 14.740 1.190 ;
        RECT  10.630 1.620 14.480 1.860 ;
        RECT  12.170 0.940 14.340 1.180 ;
        RECT  13.650 2.610 14.050 3.010 ;
        RECT  11.190 2.620 13.650 2.860 ;
        RECT  11.770 0.780 12.170 1.180 ;
        RECT  11.770 3.940 12.010 4.320 ;
        RECT  10.880 4.080 11.770 4.320 ;
        RECT  11.430 3.300 11.670 3.700 ;
        RECT  11.150 2.620 11.190 3.020 ;
        RECT  10.910 2.620 11.150 3.660 ;
        RECT  5.900 3.420 10.910 3.660 ;
        RECT  10.640 3.940 10.880 4.320 ;
        RECT  2.980 3.940 10.640 4.180 ;
        RECT  10.390 1.160 10.630 3.140 ;
        RECT  9.730 1.160 10.390 1.570 ;
        RECT  9.230 2.900 10.390 3.140 ;
        RECT  9.870 2.180 10.110 2.580 ;
        RECT  8.490 2.180 9.870 2.420 ;
        RECT  9.490 0.680 9.730 1.570 ;
        RECT  9.140 0.680 9.490 0.920 ;
        RECT  8.830 2.840 9.230 3.140 ;
        RECT  8.330 2.180 8.490 3.080 ;
        RECT  8.090 0.980 8.330 3.080 ;
        RECT  7.720 0.980 8.090 1.220 ;
        RECT  7.520 2.260 8.090 2.500 ;
        RECT  6.420 1.460 7.580 1.700 ;
        RECT  7.120 2.100 7.520 2.500 ;
        RECT  6.180 0.800 6.420 3.140 ;
        RECT  5.500 0.800 6.180 1.040 ;
        RECT  5.660 1.660 5.900 3.660 ;
        RECT  5.440 1.660 5.660 2.060 ;
        RECT  1.120 3.420 5.660 3.660 ;
        RECT  5.140 2.740 5.380 3.140 ;
        RECT  4.740 0.710 5.140 1.110 ;
        RECT  2.250 2.900 5.140 3.140 ;
        RECT  2.460 0.870 4.740 1.110 ;
        RECT  4.120 2.180 4.360 2.620 ;
        RECT  3.110 2.380 4.120 2.620 ;
        RECT  2.870 1.470 3.110 2.620 ;
        RECT  2.580 3.940 2.980 4.340 ;
        RECT  1.700 1.470 2.870 1.710 ;
        RECT  2.220 0.730 2.460 1.110 ;
        RECT  1.750 0.730 2.220 0.970 ;
        RECT  1.700 2.830 1.910 3.070 ;
        RECT  1.460 1.470 1.700 3.070 ;
        RECT  0.880 1.280 1.120 3.900 ;
        RECT  0.570 1.280 0.880 1.520 ;
        RECT  0.170 3.500 0.880 3.900 ;
        RECT  0.170 1.120 0.570 1.520 ;
    END
END EDFFX4

MACRO EDFFX2
    CLASS CORE ;
    FOREIGN EDFFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ EDFFXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.590 2.880 16.610 3.280 ;
        RECT  16.610 2.880 16.700 3.630 ;
        RECT  16.700 2.880 16.750 3.770 ;
        RECT  16.590 1.280 16.750 1.680 ;
        RECT  16.750 1.280 16.960 3.770 ;
        RECT  16.960 1.280 16.990 3.630 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.280 1.340 15.520 3.280 ;
        RECT  15.520 2.950 15.640 3.210 ;
        RECT  15.640 2.960 15.680 3.200 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 3.930 1.870 4.340 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.080 1.970 4.480 2.380 ;
        RECT  4.480 2.140 4.740 2.380 ;
        RECT  4.740 2.140 4.820 2.640 ;
        RECT  4.820 2.140 4.980 2.650 ;
        RECT  4.980 2.390 5.080 2.650 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.690 2.090 0.860 2.640 ;
        RECT  0.860 2.090 0.930 2.650 ;
        RECT  0.930 2.390 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.840 5.440 ;
        RECT  0.840 3.170 1.160 5.440 ;
        RECT  1.160 3.170 1.290 3.580 ;
        RECT  1.290 3.180 1.330 3.580 ;
        RECT  1.160 4.640 3.730 5.440 ;
        RECT  3.730 4.480 4.130 5.440 ;
        RECT  4.130 4.640 7.280 5.440 ;
        RECT  7.280 4.480 7.680 5.440 ;
        RECT  7.680 4.640 8.980 5.440 ;
        RECT  8.980 4.480 9.960 5.440 ;
        RECT  9.960 4.640 12.330 5.440 ;
        RECT  12.330 4.480 13.870 5.440 ;
        RECT  13.870 4.640 16.060 5.440 ;
        RECT  16.060 4.110 16.300 5.440 ;
        RECT  16.300 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.950 0.400 ;
        RECT  0.950 -0.400 1.350 0.560 ;
        RECT  1.350 -0.400 3.130 0.400 ;
        RECT  3.130 -0.400 3.530 0.560 ;
        RECT  3.530 -0.400 6.740 0.400 ;
        RECT  6.740 -0.400 6.750 1.130 ;
        RECT  6.750 -0.400 7.150 1.330 ;
        RECT  7.150 -0.400 7.160 1.130 ;
        RECT  7.160 -0.400 9.500 0.400 ;
        RECT  9.500 -0.400 9.900 0.560 ;
        RECT  9.900 -0.400 12.090 0.400 ;
        RECT  12.090 -0.400 12.490 0.560 ;
        RECT  12.490 -0.400 13.720 0.400 ;
        RECT  13.720 -0.400 14.120 0.560 ;
        RECT  14.120 -0.400 15.870 0.400 ;
        RECT  15.870 -0.400 16.270 0.560 ;
        RECT  16.270 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.310 2.190 16.510 2.600 ;
        RECT  16.070 2.190 16.310 3.830 ;
        RECT  15.000 3.590 16.070 3.830 ;
        RECT  14.760 0.680 15.000 4.020 ;
        RECT  14.550 0.680 14.760 0.920 ;
        RECT  14.550 3.620 14.760 4.020 ;
        RECT  13.650 3.620 14.550 3.860 ;
        RECT  13.930 2.220 14.410 2.620 ;
        RECT  13.690 1.320 13.930 2.980 ;
        RECT  13.010 1.320 13.690 1.560 ;
        RECT  13.230 2.740 13.690 2.980 ;
        RECT  13.250 3.620 13.650 4.180 ;
        RECT  12.930 1.860 13.330 2.260 ;
        RECT  2.690 3.940 13.250 4.180 ;
        RECT  12.970 2.740 13.230 3.140 ;
        RECT  12.610 1.160 13.010 1.560 ;
        RECT  12.730 2.740 12.970 3.500 ;
        RECT  12.440 2.010 12.930 2.250 ;
        RECT  11.310 3.260 12.730 3.500 ;
        RECT  11.190 1.230 12.610 1.470 ;
        RECT  12.200 2.010 12.440 2.670 ;
        RECT  11.030 2.430 12.200 2.670 ;
        RECT  11.000 1.750 11.400 2.150 ;
        RECT  10.910 3.260 11.310 3.660 ;
        RECT  10.790 1.070 11.190 1.470 ;
        RECT  10.630 2.430 11.030 2.870 ;
        RECT  10.000 1.750 11.000 1.990 ;
        RECT  10.390 2.430 10.630 3.660 ;
        RECT  5.950 3.420 10.390 3.660 ;
        RECT  9.990 1.690 10.000 1.990 ;
        RECT  9.750 1.690 9.990 3.140 ;
        RECT  9.080 1.690 9.750 1.930 ;
        RECT  8.990 2.900 9.750 3.140 ;
        RECT  9.280 2.220 9.470 2.620 ;
        RECT  8.560 2.210 9.280 2.620 ;
        RECT  8.840 0.670 9.080 1.930 ;
        RECT  8.390 0.670 8.840 0.910 ;
        RECT  8.320 1.750 8.560 3.080 ;
        RECT  8.050 1.750 8.320 1.990 ;
        RECT  8.150 2.840 8.320 3.080 ;
        RECT  7.810 0.970 8.050 1.990 ;
        RECT  6.470 2.270 8.030 2.510 ;
        RECT  6.760 1.750 7.810 1.990 ;
        RECT  6.230 1.000 6.470 3.140 ;
        RECT  5.350 1.000 6.230 1.240 ;
        RECT  5.710 1.600 5.950 3.660 ;
        RECT  5.010 1.600 5.710 1.840 ;
        RECT  5.190 3.200 5.430 3.600 ;
        RECT  2.840 3.360 5.190 3.600 ;
        RECT  4.770 1.380 5.010 1.840 ;
        RECT  2.460 0.860 4.870 1.100 ;
        RECT  0.570 1.380 4.770 1.620 ;
        RECT  3.800 2.770 4.460 3.010 ;
        RECT  3.560 1.900 3.800 3.010 ;
        RECT  2.090 1.900 3.560 2.140 ;
        RECT  2.440 3.260 2.840 3.660 ;
        RECT  2.220 0.710 2.460 1.100 ;
        RECT  1.780 0.710 2.220 0.950 ;
        RECT  1.850 1.900 2.090 3.580 ;
        RECT  1.650 1.900 1.850 2.140 ;
        RECT  1.690 3.180 1.850 3.580 ;
        RECT  0.410 1.290 0.570 1.690 ;
        RECT  0.410 3.340 0.570 3.740 ;
        RECT  0.170 1.290 0.410 3.740 ;
    END
END EDFFX2

MACRO EDFFX1
    CLASS CORE ;
    FOREIGN EDFFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ EDFFXL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.600 1.410 14.610 1.830 ;
        RECT  14.610 1.320 14.720 1.830 ;
        RECT  14.610 2.980 14.730 3.380 ;
        RECT  14.720 1.320 14.730 2.090 ;
        RECT  14.730 1.320 14.970 3.380 ;
        RECT  14.970 1.320 14.980 2.090 ;
        RECT  14.970 2.980 15.010 3.380 ;
        RECT  14.980 1.320 15.010 1.840 ;
        RECT  15.010 1.410 15.020 1.840 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.150 3.830 13.310 4.230 ;
        RECT  12.950 0.690 13.350 1.100 ;
        RECT  13.310 3.530 13.400 4.230 ;
        RECT  13.400 3.510 13.550 4.230 ;
        RECT  13.550 3.510 13.660 3.770 ;
        RECT  13.660 3.510 14.090 3.750 ;
        RECT  13.350 0.860 14.090 1.100 ;
        RECT  14.090 0.860 14.330 3.750 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 3.960 2.000 4.360 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.080 2.050 4.480 2.450 ;
        RECT  4.480 2.210 4.740 2.450 ;
        RECT  4.740 2.210 4.820 2.640 ;
        RECT  4.820 2.210 4.980 2.650 ;
        RECT  4.980 2.390 5.080 2.650 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.690 2.400 0.860 3.000 ;
        RECT  0.860 2.390 0.930 3.000 ;
        RECT  0.930 2.390 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.780 5.440 ;
        RECT  0.780 4.480 1.180 5.440 ;
        RECT  1.180 4.640 3.730 5.440 ;
        RECT  3.730 4.480 4.130 5.440 ;
        RECT  4.130 4.640 7.280 5.440 ;
        RECT  7.280 4.480 7.680 5.440 ;
        RECT  7.680 4.640 8.880 5.440 ;
        RECT  8.880 4.480 9.860 5.440 ;
        RECT  9.860 4.640 12.330 5.440 ;
        RECT  12.330 4.480 12.730 5.440 ;
        RECT  12.730 4.640 13.880 5.440 ;
        RECT  13.880 4.480 14.280 5.440 ;
        RECT  14.280 4.640 15.180 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.950 0.400 ;
        RECT  0.950 -0.400 1.350 0.560 ;
        RECT  1.350 -0.400 3.400 0.400 ;
        RECT  3.400 -0.400 3.800 0.560 ;
        RECT  3.800 -0.400 6.960 0.400 ;
        RECT  6.960 -0.400 7.360 1.280 ;
        RECT  7.360 -0.400 9.570 0.400 ;
        RECT  9.570 -0.400 9.580 0.800 ;
        RECT  9.580 -0.400 9.980 1.000 ;
        RECT  9.980 -0.400 9.990 0.800 ;
        RECT  9.990 -0.400 12.130 0.400 ;
        RECT  12.130 -0.400 12.530 0.560 ;
        RECT  12.530 -0.400 13.750 0.400 ;
        RECT  13.750 -0.400 14.150 0.560 ;
        RECT  14.150 -0.400 15.180 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  13.570 1.550 13.810 3.010 ;
        RECT  13.410 1.550 13.570 1.790 ;
        RECT  13.550 2.770 13.570 3.010 ;
        RECT  13.150 2.770 13.550 3.170 ;
        RECT  13.010 1.390 13.410 1.790 ;
        RECT  12.010 2.930 13.150 3.170 ;
        RECT  12.590 2.070 12.990 2.470 ;
        RECT  11.310 2.150 12.590 2.390 ;
        RECT  11.770 2.930 12.010 4.330 ;
        RECT  11.610 3.930 11.770 4.330 ;
        RECT  3.090 3.940 11.610 4.180 ;
        RECT  10.590 0.760 11.590 1.000 ;
        RECT  11.180 1.440 11.310 3.660 ;
        RECT  11.070 1.280 11.180 3.660 ;
        RECT  10.940 1.280 11.070 1.680 ;
        RECT  10.890 3.260 11.070 3.660 ;
        RECT  10.590 2.580 10.790 2.980 ;
        RECT  10.350 0.760 10.590 3.660 ;
        RECT  5.950 3.420 10.350 3.660 ;
        RECT  9.830 1.560 10.070 3.140 ;
        RECT  9.160 1.560 9.830 1.800 ;
        RECT  8.990 2.900 9.830 3.140 ;
        RECT  8.550 2.330 9.550 2.570 ;
        RECT  8.920 0.670 9.160 1.800 ;
        RECT  8.680 0.670 8.920 0.910 ;
        RECT  8.470 2.330 8.550 3.060 ;
        RECT  8.240 1.550 8.470 3.060 ;
        RECT  8.230 0.870 8.240 3.060 ;
        RECT  7.840 0.870 8.230 1.790 ;
        RECT  8.150 2.820 8.230 3.060 ;
        RECT  7.710 2.100 7.950 2.530 ;
        RECT  6.990 1.550 7.840 1.790 ;
        RECT  6.470 2.290 7.710 2.530 ;
        RECT  6.750 1.550 6.990 1.950 ;
        RECT  6.230 1.070 6.470 3.140 ;
        RECT  6.020 1.070 6.230 1.310 ;
        RECT  5.620 0.910 6.020 1.310 ;
        RECT  5.710 1.620 5.950 3.660 ;
        RECT  5.010 1.620 5.710 1.860 ;
        RECT  5.190 3.200 5.430 3.660 ;
        RECT  2.390 3.420 5.190 3.660 ;
        RECT  2.460 0.870 5.140 1.110 ;
        RECT  4.770 1.380 5.010 1.860 ;
        RECT  0.570 1.380 4.770 1.620 ;
        RECT  3.220 2.850 4.460 3.090 ;
        RECT  2.980 2.060 3.220 3.090 ;
        RECT  2.700 3.940 3.090 4.230 ;
        RECT  2.820 2.060 2.980 2.460 ;
        RECT  2.060 2.220 2.820 2.460 ;
        RECT  2.690 3.990 2.700 4.230 ;
        RECT  2.060 0.860 2.460 1.110 ;
        RECT  2.050 2.040 2.060 2.460 ;
        RECT  1.960 1.900 2.050 2.460 ;
        RECT  1.960 3.180 2.050 3.580 ;
        RECT  1.720 1.900 1.960 3.580 ;
        RECT  1.650 1.900 1.720 2.140 ;
        RECT  1.650 3.180 1.720 3.580 ;
        RECT  0.410 1.380 0.570 1.790 ;
        RECT  0.410 3.340 0.570 3.740 ;
        RECT  0.250 1.380 0.410 3.740 ;
        RECT  0.170 1.390 0.250 3.740 ;
    END
END EDFFX1

MACRO DLY4X1
    CLASS CORE ;
    FOREIGN DLY4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.050 3.010 4.170 3.410 ;
        RECT  4.160 2.390 4.170 2.650 ;
        RECT  4.050 1.360 4.170 1.960 ;
        RECT  4.170 1.360 4.410 3.410 ;
        RECT  4.410 2.390 4.420 2.650 ;
        RECT  4.410 3.010 4.450 3.410 ;
        RECT  4.410 1.360 4.450 1.960 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.470 2.240 0.860 2.640 ;
        RECT  0.860 2.240 0.870 2.650 ;
        RECT  0.870 2.390 1.120 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.930 5.440 ;
        RECT  0.930 4.480 1.330 5.440 ;
        RECT  1.330 4.640 3.230 5.440 ;
        RECT  3.230 4.480 3.630 5.440 ;
        RECT  3.630 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.920 0.400 ;
        RECT  0.920 -0.400 1.320 0.560 ;
        RECT  1.320 -0.400 3.230 0.400 ;
        RECT  3.230 -0.400 3.630 0.560 ;
        RECT  3.630 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.640 2.220 3.800 2.620 ;
        RECT  3.400 0.860 3.640 3.860 ;
        RECT  2.210 0.860 3.400 1.100 ;
        RECT  2.210 3.620 3.400 3.860 ;
        RECT  2.770 2.160 2.930 2.560 ;
        RECT  2.530 1.390 2.770 3.210 ;
        RECT  2.250 1.390 2.530 1.790 ;
        RECT  2.250 2.810 2.530 3.210 ;
        RECT  1.810 0.730 2.210 1.100 ;
        RECT  1.810 3.620 2.210 4.020 ;
        RECT  1.720 2.060 1.880 2.540 ;
        RECT  1.480 1.550 1.720 3.170 ;
        RECT  0.570 1.550 1.480 1.790 ;
        RECT  0.570 2.930 1.480 3.170 ;
        RECT  0.170 1.390 0.570 1.790 ;
        RECT  0.170 2.930 0.570 3.330 ;
    END
END DLY4X1

MACRO DLY3X1
    CLASS CORE ;
    FOREIGN DLY3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.050 3.010 4.170 3.410 ;
        RECT  4.160 2.390 4.170 2.650 ;
        RECT  4.050 1.360 4.170 1.960 ;
        RECT  4.170 1.360 4.410 3.410 ;
        RECT  4.410 2.390 4.420 2.650 ;
        RECT  4.410 3.010 4.450 3.410 ;
        RECT  4.410 1.360 4.450 1.960 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.470 2.240 0.860 2.640 ;
        RECT  0.860 2.240 0.870 2.650 ;
        RECT  0.870 2.390 1.120 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.010 5.440 ;
        RECT  1.010 4.480 1.410 5.440 ;
        RECT  1.410 4.640 3.230 5.440 ;
        RECT  3.230 4.480 3.630 5.440 ;
        RECT  3.630 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        RECT  0.980 -0.400 1.380 0.560 ;
        RECT  1.380 -0.400 3.230 0.400 ;
        RECT  3.230 -0.400 3.630 0.560 ;
        RECT  3.630 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.640 2.220 3.800 2.620 ;
        RECT  3.400 0.860 3.640 3.860 ;
        RECT  2.390 0.860 3.400 1.100 ;
        RECT  2.390 3.620 3.400 3.860 ;
        RECT  2.770 2.160 2.930 2.560 ;
        RECT  2.530 1.390 2.770 3.210 ;
        RECT  2.250 1.390 2.530 1.790 ;
        RECT  2.250 2.810 2.530 3.210 ;
        RECT  1.990 0.730 2.390 1.100 ;
        RECT  1.990 3.620 2.390 4.020 ;
        RECT  1.720 2.060 1.980 2.540 ;
        RECT  1.480 1.550 1.720 3.170 ;
        RECT  0.570 1.550 1.480 1.790 ;
        RECT  0.570 2.930 1.480 3.170 ;
        RECT  0.170 1.390 0.570 1.790 ;
        RECT  0.170 2.930 0.570 3.330 ;
    END
END DLY3X1

MACRO DLY2X1
    CLASS CORE ;
    FOREIGN DLY2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.050 3.010 4.170 3.410 ;
        RECT  4.160 2.390 4.170 2.650 ;
        RECT  4.050 1.360 4.170 1.960 ;
        RECT  4.170 1.360 4.410 3.410 ;
        RECT  4.410 2.390 4.420 2.650 ;
        RECT  4.410 3.010 4.450 3.410 ;
        RECT  4.410 1.360 4.450 1.960 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.470 2.240 0.860 2.640 ;
        RECT  0.860 2.240 0.870 2.650 ;
        RECT  0.870 2.390 1.120 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.070 5.440 ;
        RECT  1.070 4.480 1.470 5.440 ;
        RECT  1.470 4.640 3.230 5.440 ;
        RECT  3.230 4.480 3.630 5.440 ;
        RECT  3.630 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        RECT  0.980 -0.400 1.380 0.560 ;
        RECT  1.380 -0.400 3.230 0.400 ;
        RECT  3.230 -0.400 3.630 0.560 ;
        RECT  3.630 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.640 2.220 3.800 2.620 ;
        RECT  3.400 0.860 3.640 3.790 ;
        RECT  2.570 0.860 3.400 1.100 ;
        RECT  2.570 3.550 3.400 3.790 ;
        RECT  2.770 2.160 2.930 2.560 ;
        RECT  2.530 1.390 2.770 3.210 ;
        RECT  2.170 0.730 2.570 1.100 ;
        RECT  2.170 3.550 2.570 3.950 ;
        RECT  2.150 1.390 2.530 1.790 ;
        RECT  2.150 2.810 2.530 3.210 ;
        RECT  1.720 2.060 1.970 2.540 ;
        RECT  1.480 1.550 1.720 3.170 ;
        RECT  0.570 1.550 1.480 1.790 ;
        RECT  0.570 2.930 1.480 3.170 ;
        RECT  0.170 1.390 0.570 1.790 ;
        RECT  0.170 2.930 0.570 3.330 ;
    END
END DLY2X1

MACRO DLY1X1
    CLASS CORE ;
    FOREIGN DLY1X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.050 3.010 4.170 3.410 ;
        RECT  4.160 2.390 4.170 2.650 ;
        RECT  4.050 1.360 4.170 1.960 ;
        RECT  4.170 1.360 4.410 3.410 ;
        RECT  4.410 2.390 4.420 2.650 ;
        RECT  4.410 3.010 4.450 3.410 ;
        RECT  4.410 1.360 4.450 1.960 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.470 2.240 0.860 2.640 ;
        RECT  0.860 2.240 0.870 2.650 ;
        RECT  0.870 2.390 1.120 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.070 5.440 ;
        RECT  1.070 4.480 1.470 5.440 ;
        RECT  1.470 4.640 3.230 5.440 ;
        RECT  3.230 4.480 3.630 5.440 ;
        RECT  3.630 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.020 0.400 ;
        RECT  1.020 -0.400 1.420 0.560 ;
        RECT  1.420 -0.400 3.230 0.400 ;
        RECT  3.230 -0.400 3.630 0.560 ;
        RECT  3.630 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.640 2.220 3.800 2.620 ;
        RECT  3.400 0.860 3.640 3.790 ;
        RECT  2.660 0.860 3.400 1.100 ;
        RECT  2.660 3.550 3.400 3.790 ;
        RECT  2.770 2.160 2.930 2.560 ;
        RECT  2.530 1.550 2.770 3.050 ;
        RECT  2.260 0.730 2.660 1.100 ;
        RECT  2.260 3.550 2.660 3.950 ;
        RECT  2.400 1.550 2.530 1.790 ;
        RECT  2.400 2.810 2.530 3.050 ;
        RECT  2.000 1.390 2.400 1.790 ;
        RECT  2.000 2.810 2.400 3.210 ;
        RECT  1.720 2.100 1.970 2.500 ;
        RECT  1.480 1.550 1.720 3.170 ;
        RECT  0.570 1.550 1.480 1.790 ;
        RECT  0.570 2.930 1.480 3.170 ;
        RECT  0.170 1.390 0.570 1.790 ;
        RECT  0.170 2.930 0.570 3.330 ;
    END
END DLY1X1

MACRO DFFTRXL
    CLASS CORE ;
    FOREIGN DFFTRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.530 1.780 2.090 ;
        RECT  1.780 1.530 1.920 1.930 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.300 1.390 11.390 2.070 ;
        RECT  11.390 1.390 11.540 3.240 ;
        RECT  11.540 1.830 11.630 3.240 ;
        RECT  11.630 1.830 11.680 2.090 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.890 3.520 10.100 3.990 ;
        RECT  10.100 3.510 10.310 3.990 ;
        RECT  10.310 3.510 10.360 3.770 ;
        RECT  9.900 0.720 10.370 1.100 ;
        RECT  10.360 3.520 10.820 3.760 ;
        RECT  10.370 0.860 10.820 1.100 ;
        RECT  10.820 0.860 11.060 3.760 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.110 2.250 2.620 2.660 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.690 2.070 0.860 2.470 ;
        RECT  0.860 2.070 1.110 2.650 ;
        RECT  1.110 2.390 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.040 5.440 ;
        RECT  1.040 4.480 2.020 5.440 ;
        RECT  2.020 4.640 4.820 5.440 ;
        RECT  4.820 4.480 5.220 5.440 ;
        RECT  5.220 4.640 6.690 5.440 ;
        RECT  6.690 3.670 6.700 5.440 ;
        RECT  6.700 3.470 7.100 5.440 ;
        RECT  7.100 3.670 7.110 5.440 ;
        RECT  7.110 4.640 9.140 5.440 ;
        RECT  9.140 3.790 9.150 5.440 ;
        RECT  9.150 3.590 9.550 5.440 ;
        RECT  9.550 3.790 9.560 5.440 ;
        RECT  9.560 4.640 10.700 5.440 ;
        RECT  10.700 4.480 11.100 5.440 ;
        RECT  11.100 4.640 11.880 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.140 0.400 ;
        RECT  1.140 -0.400 1.540 0.560 ;
        RECT  1.540 -0.400 4.370 0.400 ;
        RECT  4.370 -0.400 4.380 1.320 ;
        RECT  4.380 -0.400 4.780 1.520 ;
        RECT  4.780 -0.400 4.790 1.320 ;
        RECT  4.790 -0.400 6.530 0.400 ;
        RECT  6.530 -0.400 6.540 0.950 ;
        RECT  6.540 -0.400 6.940 1.150 ;
        RECT  6.940 -0.400 6.950 0.950 ;
        RECT  6.950 -0.400 9.090 0.400 ;
        RECT  9.090 -0.400 9.490 0.560 ;
        RECT  9.490 -0.400 11.110 0.400 ;
        RECT  11.110 -0.400 11.510 0.560 ;
        RECT  11.510 -0.400 11.880 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.300 1.380 10.540 3.160 ;
        RECT  9.970 1.380 10.300 1.780 ;
        RECT  9.970 2.760 10.300 3.160 ;
        RECT  9.100 1.540 9.970 1.780 ;
        RECT  9.690 2.060 9.900 2.460 ;
        RECT  9.450 2.060 9.690 2.780 ;
        RECT  8.490 2.540 9.450 2.780 ;
        RECT  8.860 1.540 9.100 2.260 ;
        RECT  8.250 1.220 8.490 3.970 ;
        RECT  8.140 1.220 8.250 1.460 ;
        RECT  8.040 3.570 8.250 3.970 ;
        RECT  7.900 1.060 8.140 1.460 ;
        RECT  7.620 1.890 7.970 2.290 ;
        RECT  7.380 1.430 7.620 2.970 ;
        RECT  6.260 1.430 7.380 1.670 ;
        RECT  6.660 2.730 7.380 2.970 ;
        RECT  5.690 1.950 7.090 2.350 ;
        RECT  6.260 2.730 6.660 3.130 ;
        RECT  4.060 3.940 6.420 4.180 ;
        RECT  5.980 0.670 6.260 1.670 ;
        RECT  5.060 0.670 5.980 0.910 ;
        RECT  5.450 1.370 5.690 3.050 ;
        RECT  5.260 1.370 5.450 1.770 ;
        RECT  4.450 2.810 5.450 3.050 ;
        RECT  4.980 2.050 5.170 2.460 ;
        RECT  4.740 1.990 4.980 2.460 ;
        RECT  3.880 1.990 4.740 2.230 ;
        RECT  4.210 2.510 4.450 3.050 ;
        RECT  3.660 3.940 4.060 4.370 ;
        RECT  3.640 1.010 3.880 3.110 ;
        RECT  3.360 3.940 3.660 4.180 ;
        RECT  3.020 1.010 3.640 1.250 ;
        RECT  3.120 1.530 3.360 4.180 ;
        RECT  2.720 1.530 3.120 1.930 ;
        RECT  0.490 3.940 3.120 4.180 ;
        RECT  2.600 2.930 2.840 3.660 ;
        RECT  2.690 1.530 2.720 1.770 ;
        RECT  2.450 1.000 2.690 1.770 ;
        RECT  1.650 2.930 2.600 3.170 ;
        RECT  0.570 1.000 2.450 1.240 ;
        RECT  0.410 1.000 0.570 1.520 ;
        RECT  0.410 2.750 0.490 4.180 ;
        RECT  0.250 1.000 0.410 4.180 ;
        RECT  0.170 1.000 0.250 3.150 ;
    END
END DFFTRXL

MACRO DFFTRX4
    CLASS CORE ;
    FOREIGN DFFTRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFTRXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.310 1.700 1.320 2.100 ;
        RECT  1.320 1.700 1.720 2.110 ;
        RECT  1.720 1.700 1.870 2.100 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.290 1.260 15.690 3.150 ;
        RECT  15.690 1.260 15.730 2.660 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.750 2.810 13.950 3.210 ;
        RECT  13.950 1.260 13.970 3.210 ;
        RECT  13.970 1.260 14.350 3.220 ;
        RECT  14.350 1.820 14.410 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.140 2.250 2.320 2.650 ;
        RECT  2.320 2.240 2.580 2.660 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.150 0.920 2.660 ;
        RECT  0.920 2.380 1.210 2.660 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.030 5.440 ;
        RECT  1.030 4.480 1.430 5.440 ;
        RECT  1.430 4.640 5.340 5.440 ;
        RECT  5.340 4.480 5.740 5.440 ;
        RECT  5.740 4.640 6.630 5.440 ;
        RECT  6.630 4.480 7.030 5.440 ;
        RECT  7.030 4.640 9.060 5.440 ;
        RECT  9.060 3.730 9.460 5.440 ;
        RECT  9.460 4.640 11.700 5.440 ;
        RECT  11.700 4.480 11.870 5.440 ;
        RECT  11.870 3.900 12.270 5.440 ;
        RECT  12.270 4.640 13.160 5.440 ;
        RECT  13.160 4.010 13.560 5.440 ;
        RECT  13.560 4.640 14.650 5.440 ;
        RECT  14.650 4.010 15.050 5.440 ;
        RECT  15.050 4.640 15.940 5.440 ;
        RECT  15.940 4.010 16.340 5.440 ;
        RECT  16.340 4.640 16.500 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        RECT  0.990 -0.400 1.390 0.560 ;
        RECT  1.390 -0.400 4.090 0.400 ;
        RECT  4.090 -0.400 4.100 1.240 ;
        RECT  4.100 -0.400 4.500 1.440 ;
        RECT  4.500 -0.400 4.510 1.240 ;
        RECT  4.510 -0.400 6.760 0.400 ;
        RECT  6.760 -0.400 7.160 1.310 ;
        RECT  7.160 -0.400 9.190 0.400 ;
        RECT  9.190 -0.400 9.200 1.130 ;
        RECT  9.200 -0.400 9.600 1.330 ;
        RECT  9.600 -0.400 9.610 1.130 ;
        RECT  9.610 -0.400 11.840 0.400 ;
        RECT  11.840 -0.400 12.240 0.560 ;
        RECT  12.240 -0.400 13.360 0.400 ;
        RECT  13.360 -0.400 13.760 0.980 ;
        RECT  13.760 -0.400 14.650 0.400 ;
        RECT  14.650 -0.400 15.050 0.980 ;
        RECT  15.050 -0.400 15.940 0.400 ;
        RECT  15.940 -0.400 16.340 0.980 ;
        RECT  16.340 -0.400 16.500 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  15.970 2.180 16.210 3.730 ;
        RECT  13.510 3.490 15.970 3.730 ;
        RECT  13.270 1.380 13.510 3.730 ;
        RECT  13.040 1.380 13.270 1.620 ;
        RECT  12.440 2.910 13.270 3.310 ;
        RECT  12.640 1.220 13.040 1.620 ;
        RECT  12.630 2.110 13.030 2.510 ;
        RECT  12.400 2.110 12.630 2.350 ;
        RECT  11.560 3.070 12.440 3.310 ;
        RECT  12.160 1.370 12.400 2.350 ;
        RECT  10.820 1.370 12.160 1.610 ;
        RECT  11.320 3.070 11.560 3.720 ;
        RECT  11.260 1.890 11.420 2.130 ;
        RECT  11.080 1.890 11.260 2.810 ;
        RECT  11.020 1.890 11.080 4.360 ;
        RECT  10.840 2.570 11.020 4.360 ;
        RECT  10.050 4.120 10.840 4.360 ;
        RECT  10.760 1.210 10.820 1.610 ;
        RECT  10.560 1.210 10.760 2.330 ;
        RECT  10.520 1.210 10.560 3.460 ;
        RECT  10.420 1.210 10.520 1.610 ;
        RECT  10.320 2.090 10.520 3.460 ;
        RECT  8.300 2.090 10.320 2.330 ;
        RECT  9.810 3.210 10.050 4.360 ;
        RECT  8.820 3.210 9.810 3.450 ;
        RECT  8.580 3.210 8.820 4.080 ;
        RECT  6.340 3.840 8.580 4.080 ;
        RECT  8.300 1.060 8.380 1.460 ;
        RECT  8.280 1.060 8.300 2.330 ;
        RECT  8.060 1.060 8.280 3.560 ;
        RECT  7.980 1.060 8.060 1.460 ;
        RECT  8.040 2.090 8.060 3.560 ;
        RECT  7.880 3.160 8.040 3.560 ;
        RECT  7.400 1.590 7.640 3.050 ;
        RECT  6.400 1.590 7.400 1.830 ;
        RECT  6.160 2.810 7.400 3.050 ;
        RECT  5.550 2.110 7.160 2.510 ;
        RECT  6.240 1.030 6.400 1.830 ;
        RECT  5.940 3.780 6.340 4.180 ;
        RECT  6.160 0.670 6.240 1.830 ;
        RECT  6.000 0.670 6.160 1.430 ;
        RECT  5.430 0.670 6.000 0.910 ;
        RECT  4.580 3.940 5.940 4.180 ;
        RECT  5.310 1.360 5.550 2.910 ;
        RECT  5.260 1.360 5.310 1.600 ;
        RECT  5.030 2.670 5.310 2.910 ;
        RECT  4.860 1.200 5.260 1.600 ;
        RECT  4.650 2.670 5.030 3.070 ;
        RECT  4.610 1.880 5.010 2.280 ;
        RECT  4.270 2.660 4.650 3.080 ;
        RECT  3.610 1.960 4.610 2.200 ;
        RECT  4.340 3.940 4.580 4.370 ;
        RECT  2.780 4.130 4.340 4.370 ;
        RECT  3.970 2.670 4.270 3.070 ;
        RECT  3.370 0.960 3.610 3.690 ;
        RECT  2.760 0.960 3.370 1.200 ;
        RECT  3.270 3.450 3.370 3.690 ;
        RECT  3.030 3.450 3.270 3.850 ;
        RECT  2.910 1.670 3.090 3.170 ;
        RECT  2.850 1.510 2.910 3.170 ;
        RECT  2.510 1.510 2.850 1.910 ;
        RECT  2.780 2.930 2.850 3.170 ;
        RECT  2.540 2.930 2.780 4.370 ;
        RECT  2.480 1.510 2.510 1.750 ;
        RECT  2.240 1.190 2.480 1.750 ;
        RECT  2.050 3.030 2.290 4.300 ;
        RECT  0.570 1.190 2.240 1.430 ;
        RECT  1.580 3.030 2.050 3.270 ;
        RECT  0.400 1.030 0.570 1.430 ;
        RECT  0.400 3.030 0.570 4.010 ;
        RECT  0.170 1.030 0.400 4.010 ;
        RECT  0.160 1.110 0.170 3.990 ;
    END
END DFFTRX4

MACRO DFFTRX2
    CLASS CORE ;
    FOREIGN DFFTRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFTRXL ;
    SIZE 14.520 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.610 2.090 ;
        RECT  1.610 1.710 2.010 2.110 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.400 1.270 13.510 1.530 ;
        RECT  13.510 1.260 13.950 1.530 ;
        RECT  13.950 3.140 14.110 4.120 ;
        RECT  13.950 1.010 14.110 1.530 ;
        RECT  14.110 1.010 14.350 4.120 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.430 0.860 12.510 1.260 ;
        RECT  12.510 0.860 12.750 3.160 ;
        RECT  12.750 0.860 12.830 1.280 ;
        RECT  12.750 1.830 13.000 2.090 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 2.390 2.370 2.650 ;
        RECT  2.370 2.390 2.440 2.790 ;
        RECT  2.440 2.400 2.770 2.790 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.740 2.200 1.120 2.670 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.310 5.440 ;
        RECT  1.310 4.480 1.710 5.440 ;
        RECT  1.710 4.640 4.820 5.440 ;
        RECT  4.820 4.480 5.220 5.440 ;
        RECT  5.220 4.640 6.920 5.440 ;
        RECT  6.920 4.480 7.320 5.440 ;
        RECT  7.320 4.640 9.470 5.440 ;
        RECT  9.470 4.480 9.870 5.440 ;
        RECT  9.870 4.640 13.180 5.440 ;
        RECT  13.180 4.280 13.190 5.440 ;
        RECT  13.190 4.080 13.590 5.440 ;
        RECT  13.590 4.280 13.600 5.440 ;
        RECT  13.600 4.640 14.520 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.020 0.400 ;
        RECT  1.020 -0.400 1.260 1.480 ;
        RECT  1.260 -0.400 4.200 0.400 ;
        RECT  4.200 -0.400 4.210 0.730 ;
        RECT  4.210 -0.400 4.610 0.930 ;
        RECT  4.610 -0.400 4.620 0.730 ;
        RECT  4.620 -0.400 6.430 0.400 ;
        RECT  6.430 -0.400 6.440 1.140 ;
        RECT  6.440 -0.400 6.840 1.260 ;
        RECT  6.840 -0.400 6.850 1.140 ;
        RECT  6.850 -0.400 8.940 0.400 ;
        RECT  8.940 -0.400 8.950 0.980 ;
        RECT  8.950 -0.400 9.350 1.100 ;
        RECT  9.350 -0.400 9.360 0.980 ;
        RECT  9.360 -0.400 10.850 0.400 ;
        RECT  10.850 -0.400 11.250 0.560 ;
        RECT  11.250 -0.400 13.180 0.400 ;
        RECT  13.180 -0.400 13.190 0.690 ;
        RECT  13.190 -0.400 13.590 0.890 ;
        RECT  13.590 -0.400 13.600 0.690 ;
        RECT  13.600 -0.400 14.520 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  13.640 2.190 13.810 2.590 ;
        RECT  13.400 2.190 13.640 3.780 ;
        RECT  12.250 3.540 13.400 3.780 ;
        RECT  12.230 3.540 12.250 4.070 ;
        RECT  12.070 1.630 12.230 4.070 ;
        RECT  11.990 1.060 12.070 4.070 ;
        RECT  11.670 1.060 11.990 1.870 ;
        RECT  11.850 3.670 11.990 4.070 ;
        RECT  11.470 2.350 11.710 3.170 ;
        RECT  11.030 1.630 11.670 1.870 ;
        RECT  10.510 2.930 11.470 3.170 ;
        RECT  10.790 1.630 11.030 2.030 ;
        RECT  10.310 1.380 10.510 3.170 ;
        RECT  10.270 1.380 10.310 3.250 ;
        RECT  10.090 1.380 10.270 1.620 ;
        RECT  10.230 2.850 10.270 3.250 ;
        RECT  9.910 2.850 10.230 3.340 ;
        RECT  9.690 1.220 10.090 1.620 ;
        RECT  9.750 1.900 9.990 2.570 ;
        RECT  8.510 3.100 9.910 3.340 ;
        RECT  7.830 1.900 9.750 2.140 ;
        RECT  8.670 1.380 9.690 1.620 ;
        RECT  8.430 1.220 8.670 1.620 ;
        RECT  7.940 2.430 8.610 2.670 ;
        RECT  8.270 3.100 8.510 3.500 ;
        RECT  7.990 1.220 8.430 1.460 ;
        RECT  7.750 1.060 7.990 1.460 ;
        RECT  7.700 2.430 7.940 3.560 ;
        RECT  7.420 1.820 7.830 2.140 ;
        RECT  7.310 3.320 7.700 3.560 ;
        RECT  7.180 1.590 7.420 3.040 ;
        RECT  7.070 3.320 7.310 4.180 ;
        RECT  6.020 1.590 7.180 1.830 ;
        RECT  6.790 2.800 7.180 3.040 ;
        RECT  4.450 3.940 7.070 4.180 ;
        RECT  5.980 2.110 6.900 2.510 ;
        RECT  6.550 2.800 6.790 3.520 ;
        RECT  6.310 3.280 6.550 3.520 ;
        RECT  5.780 0.670 6.020 1.830 ;
        RECT  5.740 2.110 5.980 3.660 ;
        RECT  5.560 0.670 5.780 1.140 ;
        RECT  5.490 2.110 5.740 2.350 ;
        RECT  5.570 3.420 5.740 3.660 ;
        RECT  4.900 0.670 5.560 0.910 ;
        RECT  5.250 1.610 5.490 2.350 ;
        RECT  5.210 2.640 5.450 3.120 ;
        RECT  4.450 1.610 5.250 1.850 ;
        RECT  3.930 2.880 5.210 3.120 ;
        RECT  4.210 1.610 4.450 2.600 ;
        RECT  4.210 3.940 4.450 4.260 ;
        RECT  3.410 4.020 4.210 4.260 ;
        RECT  3.690 1.260 3.930 3.740 ;
        RECT  3.090 1.260 3.690 1.500 ;
        RECT  3.170 1.830 3.410 4.260 ;
        RECT  2.770 1.830 3.170 2.070 ;
        RECT  2.370 4.020 3.170 4.260 ;
        RECT  2.650 3.070 2.890 3.740 ;
        RECT  2.090 3.070 2.650 3.310 ;
        RECT  2.130 3.590 2.370 4.260 ;
        RECT  0.570 3.590 2.130 3.830 ;
        RECT  1.690 2.930 2.090 3.310 ;
        RECT  0.410 1.150 0.570 1.550 ;
        RECT  0.410 3.060 0.570 3.830 ;
        RECT  0.330 1.150 0.410 3.830 ;
        RECT  0.170 1.150 0.330 3.460 ;
    END
END DFFTRX2

MACRO DFFTRX1
    CLASS CORE ;
    FOREIGN DFFTRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFTRXL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.530 1.780 2.090 ;
        RECT  1.780 1.530 1.920 1.930 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.390 1.170 11.420 2.070 ;
        RECT  11.390 2.970 11.430 3.370 ;
        RECT  11.420 1.170 11.430 2.090 ;
        RECT  11.430 1.170 11.630 3.370 ;
        RECT  11.630 1.830 11.670 3.370 ;
        RECT  11.670 1.830 11.680 2.090 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.970 3.520 10.100 4.110 ;
        RECT  9.900 0.670 10.310 1.100 ;
        RECT  10.100 3.510 10.360 4.110 ;
        RECT  10.360 3.520 10.370 4.110 ;
        RECT  10.370 3.520 10.820 3.760 ;
        RECT  10.310 0.860 10.820 1.100 ;
        RECT  10.820 0.860 11.060 3.760 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.110 2.250 2.620 2.660 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.690 2.070 0.860 2.640 ;
        RECT  0.860 2.070 0.930 2.650 ;
        RECT  0.930 2.390 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.980 5.440 ;
        RECT  0.980 4.480 1.980 5.440 ;
        RECT  1.980 4.640 4.820 5.440 ;
        RECT  4.820 4.480 5.220 5.440 ;
        RECT  5.220 4.640 6.690 5.440 ;
        RECT  6.690 3.890 6.700 5.440 ;
        RECT  6.700 3.690 7.100 5.440 ;
        RECT  7.100 3.890 7.110 5.440 ;
        RECT  7.110 4.640 9.160 5.440 ;
        RECT  9.160 4.170 9.170 5.440 ;
        RECT  9.170 3.970 9.570 5.440 ;
        RECT  9.570 4.170 9.580 5.440 ;
        RECT  9.580 4.640 10.700 5.440 ;
        RECT  10.700 4.480 11.100 5.440 ;
        RECT  11.100 4.640 11.880 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.140 0.400 ;
        RECT  1.140 -0.400 1.540 0.560 ;
        RECT  1.540 -0.400 4.370 0.400 ;
        RECT  4.370 -0.400 4.380 1.290 ;
        RECT  4.380 -0.400 4.780 1.490 ;
        RECT  4.780 -0.400 4.790 1.290 ;
        RECT  4.790 -0.400 6.530 0.400 ;
        RECT  6.530 -0.400 6.540 0.950 ;
        RECT  6.540 -0.400 6.940 1.150 ;
        RECT  6.940 -0.400 6.950 0.950 ;
        RECT  6.950 -0.400 9.090 0.400 ;
        RECT  9.090 -0.400 9.490 0.560 ;
        RECT  9.490 -0.400 10.650 0.400 ;
        RECT  10.650 -0.400 11.050 0.560 ;
        RECT  11.050 -0.400 11.880 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.300 1.380 10.540 3.160 ;
        RECT  9.970 1.380 10.300 1.780 ;
        RECT  9.970 2.760 10.300 3.160 ;
        RECT  9.100 1.540 9.970 1.780 ;
        RECT  9.690 2.060 9.900 2.460 ;
        RECT  9.450 2.060 9.690 2.780 ;
        RECT  8.490 2.540 9.450 2.780 ;
        RECT  8.860 1.540 9.100 2.260 ;
        RECT  8.250 1.220 8.490 3.970 ;
        RECT  8.140 1.220 8.250 1.460 ;
        RECT  7.980 3.570 8.250 3.970 ;
        RECT  7.900 1.060 8.140 1.460 ;
        RECT  7.620 1.890 7.970 2.290 ;
        RECT  7.380 1.430 7.620 2.970 ;
        RECT  6.260 1.430 7.380 1.670 ;
        RECT  6.660 2.730 7.380 2.970 ;
        RECT  5.690 1.950 7.090 2.350 ;
        RECT  6.260 2.730 6.660 3.130 ;
        RECT  4.060 3.940 6.420 4.180 ;
        RECT  5.980 0.670 6.260 1.670 ;
        RECT  5.060 0.670 5.980 0.910 ;
        RECT  5.450 1.370 5.690 3.050 ;
        RECT  5.260 1.370 5.450 1.770 ;
        RECT  4.450 2.810 5.450 3.050 ;
        RECT  4.980 2.050 5.170 2.460 ;
        RECT  4.740 1.990 4.980 2.460 ;
        RECT  3.880 1.990 4.740 2.230 ;
        RECT  4.210 2.510 4.450 3.050 ;
        RECT  3.660 3.940 4.060 4.370 ;
        RECT  3.640 1.020 3.880 3.110 ;
        RECT  3.360 3.940 3.660 4.180 ;
        RECT  3.020 1.020 3.640 1.260 ;
        RECT  3.120 1.530 3.360 4.180 ;
        RECT  2.720 1.530 3.120 1.930 ;
        RECT  0.570 3.940 3.120 4.180 ;
        RECT  2.600 2.930 2.840 3.660 ;
        RECT  2.690 1.530 2.720 1.770 ;
        RECT  2.450 0.930 2.690 1.770 ;
        RECT  1.650 2.930 2.600 3.170 ;
        RECT  0.570 0.930 2.450 1.170 ;
        RECT  0.410 0.930 0.570 1.330 ;
        RECT  0.410 2.930 0.570 4.180 ;
        RECT  0.330 0.930 0.410 4.180 ;
        RECT  0.170 0.930 0.330 3.330 ;
    END
END DFFTRX1

MACRO DFFSRHQXL
    CLASS CORE ;
    FOREIGN DFFSRHQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.420 4.130 6.190 4.370 ;
        RECT  6.190 3.570 6.430 4.370 ;
        RECT  6.430 3.570 7.230 3.810 ;
        RECT  7.230 3.570 7.470 4.370 ;
        RECT  7.470 4.130 9.990 4.370 ;
        RECT  9.990 3.660 10.230 4.370 ;
        RECT  10.230 3.660 10.350 3.900 ;
        RECT  10.350 3.520 10.450 3.900 ;
        RECT  10.450 3.500 10.630 3.900 ;
        RECT  10.630 2.390 10.870 3.900 ;
        RECT  10.870 2.390 11.050 2.700 ;
        RECT  11.050 2.460 11.130 2.700 ;
        RECT  14.020 2.340 14.310 2.580 ;
        RECT  14.310 2.340 14.410 2.640 ;
        RECT  10.870 3.660 14.590 3.900 ;
        RECT  14.410 2.340 14.590 2.660 ;
        RECT  14.590 2.340 14.830 3.900 ;
        RECT  14.830 2.640 15.070 3.020 ;
        RECT  15.070 2.700 15.360 3.020 ;
        RECT  15.360 2.620 15.760 3.020 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  12.910 2.390 13.400 2.630 ;
        RECT  13.400 2.390 13.660 2.650 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.110 3.600 15.510 4.000 ;
        RECT  15.510 3.600 16.040 3.840 ;
        RECT  15.100 1.270 16.040 1.540 ;
        RECT  16.040 1.270 16.080 3.840 ;
        RECT  16.080 1.280 16.280 3.840 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 1.530 1.470 1.930 ;
        RECT  1.470 1.520 1.780 2.090 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.740 2.230 0.770 2.650 ;
        RECT  0.770 2.220 1.170 2.660 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.130 5.440 ;
        RECT  1.130 4.480 1.530 5.440 ;
        RECT  1.530 4.640 3.740 5.440 ;
        RECT  3.740 4.480 4.140 5.440 ;
        RECT  4.140 4.640 6.710 5.440 ;
        RECT  6.710 4.090 6.950 5.440 ;
        RECT  6.950 4.640 10.500 5.440 ;
        RECT  10.500 4.300 10.510 5.440 ;
        RECT  10.510 4.180 10.910 5.440 ;
        RECT  10.910 4.300 10.920 5.440 ;
        RECT  10.920 4.640 12.410 5.440 ;
        RECT  12.410 4.480 12.810 5.440 ;
        RECT  12.810 4.640 13.830 5.440 ;
        RECT  13.830 4.480 14.230 5.440 ;
        RECT  14.230 4.640 15.930 5.440 ;
        RECT  15.930 4.480 16.330 5.440 ;
        RECT  16.330 4.640 16.500 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.030 0.400 ;
        RECT  1.030 -0.400 1.430 0.560 ;
        RECT  1.430 -0.400 3.610 0.400 ;
        RECT  3.610 -0.400 3.620 0.730 ;
        RECT  3.620 -0.400 4.020 0.850 ;
        RECT  4.020 -0.400 4.030 0.730 ;
        RECT  4.030 -0.400 7.300 0.400 ;
        RECT  7.300 -0.400 7.310 0.730 ;
        RECT  7.310 -0.400 7.710 0.850 ;
        RECT  7.710 -0.400 7.720 0.730 ;
        RECT  7.720 -0.400 10.040 0.400 ;
        RECT  10.040 -0.400 10.440 0.560 ;
        RECT  10.440 -0.400 13.520 0.400 ;
        RECT  13.520 -0.400 13.530 0.760 ;
        RECT  13.530 -0.400 13.930 0.880 ;
        RECT  13.930 -0.400 13.940 0.760 ;
        RECT  13.940 -0.400 16.500 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.750 0.750 16.330 0.990 ;
        RECT  15.310 1.820 15.710 2.300 ;
        RECT  13.190 1.820 15.310 2.060 ;
        RECT  14.510 0.750 14.750 1.540 ;
        RECT  14.350 1.140 14.510 1.540 ;
        RECT  14.070 2.960 14.310 3.380 ;
        RECT  12.620 2.960 14.070 3.200 ;
        RECT  12.950 1.320 13.190 2.060 ;
        RECT  11.570 0.670 13.100 0.910 ;
        RECT  12.620 1.820 12.950 2.060 ;
        RECT  12.380 1.820 12.620 3.200 ;
        RECT  12.100 1.970 12.380 2.370 ;
        RECT  11.680 1.450 11.870 1.690 ;
        RECT  11.440 1.450 11.680 3.380 ;
        RECT  11.250 0.670 11.570 1.120 ;
        RECT  10.330 1.450 11.440 1.690 ;
        RECT  11.200 2.980 11.440 3.380 ;
        RECT  11.170 0.860 11.250 1.120 ;
        RECT  9.810 0.860 11.170 1.100 ;
        RECT  10.090 1.450 10.330 2.680 ;
        RECT  9.570 0.860 9.810 3.270 ;
        RECT  9.310 3.510 9.710 3.850 ;
        RECT  9.300 0.860 9.570 1.130 ;
        RECT  8.960 3.030 9.570 3.270 ;
        RECT  7.950 3.510 9.310 3.750 ;
        RECT  8.810 0.890 9.300 1.130 ;
        RECT  9.050 1.430 9.290 2.750 ;
        RECT  8.310 1.430 9.050 1.670 ;
        RECT  8.600 2.510 9.050 2.750 ;
        RECT  7.950 1.950 8.740 2.190 ;
        RECT  8.280 2.510 8.600 3.250 ;
        RECT  8.070 1.270 8.310 1.670 ;
        RECT  8.200 2.920 8.280 3.250 ;
        RECT  7.790 1.950 7.950 3.750 ;
        RECT  7.710 1.130 7.790 3.750 ;
        RECT  7.550 1.130 7.710 2.190 ;
        RECT  6.560 2.930 7.710 3.170 ;
        RECT  6.830 1.130 7.550 1.370 ;
        RECT  7.030 1.770 7.270 2.570 ;
        RECT  5.390 1.770 7.030 2.010 ;
        RECT  6.670 1.130 6.830 1.490 ;
        RECT  6.430 0.670 6.670 1.490 ;
        RECT  5.910 2.290 6.460 2.530 ;
        RECT  6.260 0.670 6.430 0.910 ;
        RECT  5.670 2.290 5.910 3.850 ;
        RECT  3.410 3.610 5.670 3.850 ;
        RECT  5.150 1.270 5.390 3.330 ;
        RECT  5.110 1.270 5.150 1.670 ;
        RECT  3.790 3.090 5.150 3.330 ;
        RECT  4.630 2.000 4.870 2.410 ;
        RECT  3.000 2.000 4.630 2.240 ;
        RECT  3.550 2.520 3.790 3.330 ;
        RECT  3.390 2.520 3.550 2.760 ;
        RECT  3.170 3.610 3.410 4.370 ;
        RECT  2.200 4.130 3.170 4.370 ;
        RECT  2.760 1.250 3.000 3.330 ;
        RECT  2.690 1.250 2.760 1.570 ;
        RECT  2.720 3.090 2.760 3.330 ;
        RECT  2.480 3.090 2.720 3.850 ;
        RECT  2.450 1.170 2.690 1.570 ;
        RECT  2.200 1.860 2.400 2.810 ;
        RECT  2.160 1.860 2.200 4.370 ;
        RECT  1.960 2.570 2.160 4.370 ;
        RECT  0.490 3.160 1.960 3.400 ;
        RECT  0.670 1.390 1.070 1.790 ;
        RECT  0.450 1.550 0.670 1.790 ;
        RECT  0.450 3.080 0.490 3.480 ;
        RECT  0.210 1.550 0.450 3.480 ;
    END
END DFFSRHQXL

MACRO DFFSRHQX4
    CLASS CORE ;
    FOREIGN DFFSRHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSRHQXL ;
    SIZE 25.080 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.580 4.130 6.880 4.370 ;
        RECT  6.880 3.660 7.150 4.370 ;
        RECT  7.150 3.660 10.010 3.900 ;
        RECT  10.010 3.660 10.250 4.370 ;
        RECT  10.250 4.130 13.580 4.370 ;
        RECT  13.580 3.660 13.820 4.370 ;
        RECT  13.820 3.660 14.060 3.900 ;
        RECT  14.060 2.460 14.400 3.900 ;
        RECT  14.400 2.460 14.460 2.700 ;
        RECT  14.400 3.660 17.470 3.900 ;
        RECT  17.470 3.020 17.710 3.900 ;
        RECT  17.710 3.020 22.060 3.260 ;
        RECT  22.060 2.340 22.300 3.260 ;
        RECT  22.300 2.340 22.970 2.580 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  16.520 2.320 16.620 2.720 ;
        RECT  16.620 2.310 17.220 2.730 ;
        RECT  17.220 2.320 17.500 2.720 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.230 3.540 18.810 3.940 ;
        RECT  18.770 1.390 20.420 1.630 ;
        RECT  18.810 3.540 20.670 3.780 ;
        RECT  20.420 1.310 20.820 1.710 ;
        RECT  20.670 3.540 21.070 3.940 ;
        RECT  20.820 1.390 22.110 1.630 ;
        RECT  22.110 1.310 22.270 1.710 ;
        RECT  22.270 1.310 22.510 2.060 ;
        RECT  21.070 3.540 22.650 3.780 ;
        RECT  22.510 1.820 22.770 2.060 ;
        RECT  22.650 3.000 22.780 3.980 ;
        RECT  22.780 2.940 23.050 3.980 ;
        RECT  23.050 2.940 23.210 3.400 ;
        RECT  22.770 1.820 23.210 2.100 ;
        RECT  23.210 1.820 23.610 3.400 ;
        RECT  23.610 1.820 23.650 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.310 1.550 1.520 1.950 ;
        RECT  1.520 1.550 1.770 2.090 ;
        RECT  1.770 1.830 1.780 2.090 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.700 2.270 1.100 2.780 ;
        RECT  1.100 2.380 1.210 2.780 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.080 5.440 ;
        RECT  1.080 3.900 1.480 5.440 ;
        RECT  1.480 4.640 3.900 5.440 ;
        RECT  3.900 4.480 4.300 5.440 ;
        RECT  4.300 4.640 7.390 5.440 ;
        RECT  7.390 4.310 7.400 5.440 ;
        RECT  7.400 4.190 7.800 5.440 ;
        RECT  7.800 4.310 7.810 5.440 ;
        RECT  7.810 4.640 9.090 5.440 ;
        RECT  9.090 4.300 9.100 5.440 ;
        RECT  9.100 4.180 9.500 5.440 ;
        RECT  9.500 4.300 9.510 5.440 ;
        RECT  9.510 4.640 14.090 5.440 ;
        RECT  14.090 4.300 14.100 5.440 ;
        RECT  14.100 4.180 14.500 5.440 ;
        RECT  14.500 4.300 14.510 5.440 ;
        RECT  14.510 4.640 15.950 5.440 ;
        RECT  15.950 4.480 16.350 5.440 ;
        RECT  16.350 4.640 17.610 5.440 ;
        RECT  17.610 4.480 18.010 5.440 ;
        RECT  18.010 4.640 19.440 5.440 ;
        RECT  19.440 4.320 19.450 5.440 ;
        RECT  19.450 4.120 19.850 5.440 ;
        RECT  19.850 4.320 19.860 5.440 ;
        RECT  19.860 4.640 21.880 5.440 ;
        RECT  21.880 4.320 21.890 5.440 ;
        RECT  21.890 4.120 22.290 5.440 ;
        RECT  22.290 4.320 22.300 5.440 ;
        RECT  22.300 4.640 23.400 5.440 ;
        RECT  23.400 4.160 23.410 5.440 ;
        RECT  23.410 3.960 23.810 5.440 ;
        RECT  23.810 4.160 23.820 5.440 ;
        RECT  23.820 4.640 25.080 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.920 0.400 ;
        RECT  0.920 -0.400 0.930 0.740 ;
        RECT  0.930 -0.400 1.330 0.940 ;
        RECT  1.330 -0.400 1.340 0.740 ;
        RECT  1.340 -0.400 3.710 0.400 ;
        RECT  3.710 -0.400 3.950 0.930 ;
        RECT  3.950 -0.400 7.580 0.400 ;
        RECT  7.580 -0.400 7.590 0.980 ;
        RECT  7.590 -0.400 7.990 1.100 ;
        RECT  7.990 -0.400 8.000 0.980 ;
        RECT  8.000 -0.400 9.160 0.400 ;
        RECT  9.160 -0.400 9.170 1.110 ;
        RECT  9.170 -0.400 9.570 1.230 ;
        RECT  9.570 -0.400 9.580 1.110 ;
        RECT  9.580 -0.400 13.560 0.400 ;
        RECT  13.560 -0.400 13.960 0.560 ;
        RECT  13.960 -0.400 17.220 0.400 ;
        RECT  17.220 -0.400 17.620 1.320 ;
        RECT  17.620 -0.400 23.770 0.400 ;
        RECT  23.770 -0.400 24.170 0.560 ;
        RECT  24.170 -0.400 25.080 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  24.420 1.280 24.820 1.680 ;
        RECT  23.100 1.280 24.420 1.520 ;
        RECT  22.860 0.750 23.100 1.520 ;
        RECT  21.760 0.750 22.860 0.990 ;
        RECT  21.360 0.670 21.760 1.070 ;
        RECT  21.270 1.960 21.670 2.360 ;
        RECT  19.930 0.750 21.360 0.990 ;
        RECT  19.830 2.040 21.270 2.280 ;
        RECT  19.530 0.670 19.930 1.070 ;
        RECT  19.820 2.040 19.830 2.540 ;
        RECT  19.420 2.040 19.820 2.730 ;
        RECT  19.410 2.040 19.420 2.540 ;
        RECT  18.450 2.040 19.410 2.280 ;
        RECT  18.340 1.770 18.450 2.280 ;
        RECT  18.210 1.320 18.340 2.280 ;
        RECT  17.940 1.320 18.210 2.010 ;
        RECT  16.930 1.770 17.940 2.010 ;
        RECT  15.950 3.080 17.190 3.320 ;
        RECT  16.900 1.400 16.930 2.010 ;
        RECT  16.500 1.320 16.900 2.010 ;
        RECT  15.070 0.730 16.570 0.970 ;
        RECT  15.950 1.770 16.500 2.010 ;
        RECT  15.710 1.770 15.950 3.320 ;
        RECT  15.010 1.460 15.370 1.700 ;
        RECT  14.750 0.730 15.070 1.120 ;
        RECT  14.770 1.460 15.010 3.380 ;
        RECT  13.610 1.460 14.770 1.700 ;
        RECT  14.690 2.980 14.770 3.380 ;
        RECT  14.670 0.860 14.750 1.120 ;
        RECT  12.620 0.860 14.670 1.100 ;
        RECT  13.370 1.460 13.610 2.240 ;
        RECT  12.980 3.560 13.300 3.800 ;
        RECT  12.730 3.560 12.980 3.830 ;
        RECT  12.450 2.880 12.950 3.280 ;
        RECT  10.810 3.590 12.730 3.830 ;
        RECT  12.450 0.860 12.620 1.570 ;
        RECT  12.210 0.670 12.450 3.310 ;
        RECT  11.110 0.670 12.210 0.910 ;
        RECT  11.090 3.070 12.210 3.310 ;
        RECT  11.700 1.250 11.860 1.490 ;
        RECT  11.460 1.250 11.700 1.750 ;
        RECT  11.050 1.510 11.460 1.750 ;
        RECT  10.870 0.670 11.110 1.230 ;
        RECT  10.810 1.510 11.050 2.790 ;
        RECT  10.700 0.990 10.870 1.230 ;
        RECT  10.330 1.510 10.810 1.750 ;
        RECT  10.460 2.550 10.810 2.790 ;
        RECT  10.570 3.140 10.810 3.830 ;
        RECT  8.000 3.140 10.570 3.380 ;
        RECT  8.000 2.030 10.530 2.270 ;
        RECT  10.140 2.550 10.460 2.860 ;
        RECT  9.930 1.170 10.330 1.750 ;
        RECT  8.280 2.620 10.140 2.860 ;
        RECT  8.810 1.510 9.930 1.750 ;
        RECT  8.410 1.170 8.810 1.750 ;
        RECT  7.990 1.380 8.000 2.270 ;
        RECT  7.990 3.000 8.000 3.380 ;
        RECT  7.760 1.380 7.990 3.380 ;
        RECT  7.120 1.380 7.760 1.620 ;
        RECT  7.750 2.030 7.760 3.380 ;
        RECT  6.900 3.000 7.750 3.240 ;
        RECT  7.220 1.900 7.460 2.570 ;
        RECT  6.060 1.900 7.220 2.140 ;
        RECT  6.700 0.660 7.120 1.630 ;
        RECT  6.580 2.420 6.820 2.660 ;
        RECT  6.410 0.670 6.700 0.910 ;
        RECT  6.340 2.420 6.580 3.850 ;
        RECT  6.130 1.220 6.370 1.620 ;
        RECT  3.620 3.610 6.340 3.850 ;
        RECT  5.890 0.750 6.130 1.620 ;
        RECT  5.820 1.900 6.060 3.230 ;
        RECT  4.850 0.750 5.890 0.990 ;
        RECT  5.610 1.900 5.820 2.140 ;
        RECT  3.950 2.990 5.820 3.230 ;
        RECT  5.350 1.270 5.610 2.140 ;
        RECT  4.840 2.420 5.390 2.660 ;
        RECT  5.210 1.270 5.350 1.670 ;
        RECT  4.610 0.750 4.850 1.630 ;
        RECT  4.600 1.910 4.840 2.660 ;
        RECT  4.450 1.230 4.610 1.630 ;
        RECT  3.050 1.910 4.600 2.150 ;
        RECT  3.710 2.520 3.950 3.230 ;
        RECT  3.490 2.520 3.710 2.760 ;
        RECT  3.380 3.610 3.620 4.350 ;
        RECT  2.380 4.110 3.380 4.350 ;
        RECT  2.900 1.030 3.050 2.730 ;
        RECT  2.810 1.030 2.900 3.550 ;
        RECT  2.670 1.030 2.810 1.270 ;
        RECT  2.660 2.490 2.810 3.550 ;
        RECT  2.270 0.870 2.670 1.270 ;
        RECT  2.140 1.730 2.380 4.350 ;
        RECT  2.120 3.380 2.140 4.350 ;
        RECT  0.570 3.380 2.120 3.620 ;
        RECT  0.410 1.120 0.570 1.520 ;
        RECT  0.410 3.200 0.570 4.180 ;
        RECT  0.170 1.120 0.410 4.180 ;
    END
END DFFSRHQX4

MACRO DFFSRHQX2
    CLASS CORE ;
    FOREIGN DFFSRHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSRHQXL ;
    SIZE 21.780 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.420 4.130 6.190 4.370 ;
        RECT  6.190 3.660 6.430 4.370 ;
        RECT  6.430 3.660 9.450 3.900 ;
        RECT  9.450 3.660 9.620 4.080 ;
        RECT  9.620 3.660 9.860 4.370 ;
        RECT  9.860 4.130 13.100 4.370 ;
        RECT  13.100 3.660 13.320 4.370 ;
        RECT  13.320 2.540 13.340 4.370 ;
        RECT  13.340 2.540 13.610 3.900 ;
        RECT  13.610 2.380 13.750 3.900 ;
        RECT  13.750 2.380 14.010 2.780 ;
        RECT  13.750 3.660 14.910 3.900 ;
        RECT  14.910 3.610 15.150 3.900 ;
        RECT  15.150 3.610 17.350 3.850 ;
        RECT  17.350 3.020 17.590 3.850 ;
        RECT  17.590 3.020 18.930 3.260 ;
        RECT  18.930 2.940 19.080 3.260 ;
        RECT  19.080 2.770 19.470 3.260 ;
        RECT  19.470 2.770 19.850 3.010 ;
        RECT  19.850 2.040 20.090 3.010 ;
        RECT  20.090 2.040 20.290 2.280 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  15.950 2.310 16.550 2.730 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.440 3.540 18.840 3.940 ;
        RECT  18.630 1.390 19.030 1.760 ;
        RECT  18.840 3.540 19.460 3.780 ;
        RECT  19.460 3.500 19.910 3.780 ;
        RECT  19.910 3.500 20.540 3.790 ;
        RECT  20.540 3.000 20.570 3.980 ;
        RECT  19.030 1.520 20.570 1.760 ;
        RECT  20.570 1.520 20.810 3.980 ;
        RECT  20.810 3.000 20.940 3.980 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 1.280 1.520 2.050 ;
        RECT  1.520 1.270 1.670 2.050 ;
        RECT  1.670 1.270 1.780 1.530 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.690 2.380 1.210 2.850 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.020 5.440 ;
        RECT  1.020 4.480 1.420 5.440 ;
        RECT  1.420 4.640 3.740 5.440 ;
        RECT  3.740 4.480 4.140 5.440 ;
        RECT  4.140 4.640 6.700 5.440 ;
        RECT  6.700 4.300 6.710 5.440 ;
        RECT  6.710 4.180 7.110 5.440 ;
        RECT  7.110 4.300 7.120 5.440 ;
        RECT  7.120 4.640 8.710 5.440 ;
        RECT  8.710 4.300 8.720 5.440 ;
        RECT  8.720 4.180 9.120 5.440 ;
        RECT  9.120 4.300 9.130 5.440 ;
        RECT  9.130 4.640 13.610 5.440 ;
        RECT  13.610 4.300 13.620 5.440 ;
        RECT  13.620 4.180 14.020 5.440 ;
        RECT  14.020 4.300 14.030 5.440 ;
        RECT  14.030 4.640 15.560 5.440 ;
        RECT  15.560 4.480 15.960 5.440 ;
        RECT  15.960 4.640 17.140 5.440 ;
        RECT  17.140 4.480 17.540 5.440 ;
        RECT  17.540 4.640 19.770 5.440 ;
        RECT  19.770 4.370 19.780 5.440 ;
        RECT  19.780 4.250 20.180 5.440 ;
        RECT  20.180 4.370 20.190 5.440 ;
        RECT  20.190 4.640 21.780 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        RECT  0.990 -0.400 1.390 0.560 ;
        RECT  1.390 -0.400 3.480 0.400 ;
        RECT  3.480 -0.400 3.490 0.730 ;
        RECT  3.490 -0.400 3.890 0.850 ;
        RECT  3.890 -0.400 3.900 0.730 ;
        RECT  3.900 -0.400 7.300 0.400 ;
        RECT  7.300 -0.400 7.310 0.730 ;
        RECT  7.310 -0.400 7.710 0.850 ;
        RECT  7.710 -0.400 7.720 0.730 ;
        RECT  7.720 -0.400 8.800 0.400 ;
        RECT  8.800 -0.400 8.810 1.110 ;
        RECT  8.810 -0.400 9.210 1.230 ;
        RECT  9.210 -0.400 9.220 1.110 ;
        RECT  9.220 -0.400 13.140 0.400 ;
        RECT  13.140 -0.400 13.540 0.560 ;
        RECT  13.540 -0.400 16.900 0.400 ;
        RECT  16.900 -0.400 16.910 1.120 ;
        RECT  16.910 -0.400 17.310 1.320 ;
        RECT  17.310 -0.400 17.320 1.120 ;
        RECT  17.320 -0.400 20.650 0.400 ;
        RECT  20.650 -0.400 20.660 1.020 ;
        RECT  20.660 -0.400 21.060 1.140 ;
        RECT  21.060 -0.400 21.070 1.020 ;
        RECT  21.070 -0.400 21.780 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  18.270 0.790 19.940 1.030 ;
        RECT  17.450 2.040 19.510 2.280 ;
        RECT  18.030 0.670 18.270 1.030 ;
        RECT  17.870 0.670 18.030 0.910 ;
        RECT  17.210 1.770 17.450 2.280 ;
        RECT  16.540 1.770 17.210 2.010 ;
        RECT  15.560 3.080 16.800 3.320 ;
        RECT  16.140 1.320 16.540 2.010 ;
        RECT  14.660 0.670 16.200 0.910 ;
        RECT  15.560 1.770 16.140 2.010 ;
        RECT  15.320 1.770 15.560 3.320 ;
        RECT  14.540 1.460 14.970 1.700 ;
        RECT  14.340 0.670 14.660 1.120 ;
        RECT  14.540 3.020 14.620 3.300 ;
        RECT  14.300 1.460 14.540 3.300 ;
        RECT  14.260 0.860 14.340 1.120 ;
        RECT  13.210 1.460 14.300 1.700 ;
        RECT  14.220 3.020 14.300 3.300 ;
        RECT  12.250 0.860 14.260 1.100 ;
        RECT  12.970 1.460 13.210 2.240 ;
        RECT  10.450 3.610 12.820 3.850 ;
        RECT  12.090 2.930 12.470 3.330 ;
        RECT  12.090 0.860 12.250 1.580 ;
        RECT  11.850 0.670 12.090 3.330 ;
        RECT  10.750 0.670 11.850 0.910 ;
        RECT  10.730 3.090 11.850 3.330 ;
        RECT  11.340 1.250 11.500 1.490 ;
        RECT  11.100 1.250 11.340 1.750 ;
        RECT  10.690 1.510 11.100 1.750 ;
        RECT  10.510 0.670 10.750 1.230 ;
        RECT  10.450 1.510 10.690 2.800 ;
        RECT  10.340 0.990 10.510 1.230 ;
        RECT  9.970 1.510 10.450 1.750 ;
        RECT  9.920 2.560 10.450 2.800 ;
        RECT  10.210 3.140 10.450 3.850 ;
        RECT  7.640 3.140 10.210 3.380 ;
        RECT  7.640 2.030 10.170 2.270 ;
        RECT  9.570 1.170 9.970 1.750 ;
        RECT  9.600 2.560 9.920 2.860 ;
        RECT  7.920 2.620 9.600 2.860 ;
        RECT  8.450 1.510 9.570 1.750 ;
        RECT  8.050 1.170 8.450 1.750 ;
        RECT  7.400 1.250 7.640 3.380 ;
        RECT  6.670 1.250 7.400 1.490 ;
        RECT  6.560 2.930 7.400 3.170 ;
        RECT  6.860 1.770 7.100 2.570 ;
        RECT  5.390 1.770 6.860 2.010 ;
        RECT  6.430 0.670 6.670 1.490 ;
        RECT  5.910 2.290 6.460 2.530 ;
        RECT  6.260 0.670 6.430 0.910 ;
        RECT  5.670 2.290 5.910 3.850 ;
        RECT  3.410 3.610 5.670 3.850 ;
        RECT  5.150 1.270 5.390 3.330 ;
        RECT  5.110 1.270 5.150 1.670 ;
        RECT  3.790 3.090 5.150 3.330 ;
        RECT  4.630 2.000 4.870 2.410 ;
        RECT  3.000 2.000 4.630 2.240 ;
        RECT  3.550 2.520 3.790 3.330 ;
        RECT  3.390 2.520 3.550 2.760 ;
        RECT  3.170 3.610 3.410 4.350 ;
        RECT  2.200 4.110 3.170 4.350 ;
        RECT  2.770 1.300 3.000 2.740 ;
        RECT  2.760 1.140 2.770 2.740 ;
        RECT  2.370 1.140 2.760 1.540 ;
        RECT  2.720 2.500 2.760 2.740 ;
        RECT  2.480 2.500 2.720 3.830 ;
        RECT  2.200 1.820 2.480 2.060 ;
        RECT  1.960 1.820 2.200 4.350 ;
        RECT  0.600 3.640 1.960 3.880 ;
        RECT  0.450 3.480 0.600 3.880 ;
        RECT  0.450 1.390 0.570 1.790 ;
        RECT  0.210 1.390 0.450 3.880 ;
        RECT  0.170 1.390 0.210 1.790 ;
        RECT  0.200 3.480 0.210 3.880 ;
    END
END DFFSRHQX2

MACRO DFFSRHQX1
    CLASS CORE ;
    FOREIGN DFFSRHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSRHQXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.420 4.130 6.190 4.370 ;
        RECT  6.190 3.570 6.430 4.370 ;
        RECT  6.430 3.570 7.230 3.810 ;
        RECT  7.230 3.570 7.470 4.370 ;
        RECT  7.470 4.130 9.990 4.370 ;
        RECT  9.990 3.660 10.230 4.370 ;
        RECT  10.230 3.660 10.350 3.900 ;
        RECT  10.350 3.520 10.450 3.900 ;
        RECT  10.450 3.500 10.630 3.900 ;
        RECT  10.630 2.400 10.760 3.900 ;
        RECT  10.760 2.390 10.870 3.900 ;
        RECT  10.870 2.390 11.020 2.700 ;
        RECT  11.020 2.400 11.070 2.700 ;
        RECT  11.070 2.460 11.150 2.700 ;
        RECT  10.870 3.660 14.490 3.900 ;
        RECT  14.290 2.340 14.490 2.580 ;
        RECT  14.490 2.340 14.730 3.900 ;
        RECT  14.730 2.640 14.970 2.960 ;
        RECT  14.970 2.640 15.070 2.940 ;
        RECT  15.070 2.700 15.650 2.940 ;
        RECT  15.650 2.620 16.050 3.020 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  12.910 2.400 13.400 2.640 ;
        RECT  13.400 2.390 13.660 2.650 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.360 3.630 15.760 4.030 ;
        RECT  15.410 1.280 16.040 1.520 ;
        RECT  15.760 3.630 16.290 3.870 ;
        RECT  16.040 1.270 16.300 1.530 ;
        RECT  16.290 3.520 16.330 3.870 ;
        RECT  16.300 1.290 16.330 1.530 ;
        RECT  16.330 1.290 16.570 3.870 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.340 2.380 1.780 2.910 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.070 0.830 2.470 ;
        RECT  0.830 1.840 0.860 2.470 ;
        RECT  0.860 1.830 1.070 2.470 ;
        RECT  1.070 1.830 1.120 2.090 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.880 5.440 ;
        RECT  0.880 4.480 1.280 5.440 ;
        RECT  1.280 4.640 3.740 5.440 ;
        RECT  3.740 4.480 4.140 5.440 ;
        RECT  4.140 4.640 6.710 5.440 ;
        RECT  6.710 4.090 6.950 5.440 ;
        RECT  6.950 4.640 10.500 5.440 ;
        RECT  10.500 4.300 10.510 5.440 ;
        RECT  10.510 4.180 10.910 5.440 ;
        RECT  10.910 4.300 10.920 5.440 ;
        RECT  10.920 4.640 12.450 5.440 ;
        RECT  12.450 4.480 12.850 5.440 ;
        RECT  12.850 4.640 14.080 5.440 ;
        RECT  14.080 4.480 14.480 5.440 ;
        RECT  14.480 4.640 16.180 5.440 ;
        RECT  16.180 4.480 16.580 5.440 ;
        RECT  16.580 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.770 0.400 ;
        RECT  0.770 -0.400 1.170 0.560 ;
        RECT  1.170 -0.400 3.610 0.400 ;
        RECT  3.610 -0.400 3.620 0.730 ;
        RECT  3.620 -0.400 4.020 0.850 ;
        RECT  4.020 -0.400 4.030 0.730 ;
        RECT  4.030 -0.400 7.300 0.400 ;
        RECT  7.300 -0.400 7.310 0.730 ;
        RECT  7.310 -0.400 7.710 0.850 ;
        RECT  7.710 -0.400 7.720 0.730 ;
        RECT  7.720 -0.400 10.240 0.400 ;
        RECT  10.240 -0.400 10.640 0.560 ;
        RECT  10.640 -0.400 13.890 0.400 ;
        RECT  13.890 -0.400 14.290 1.540 ;
        RECT  14.290 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  15.050 0.750 16.630 0.990 ;
        RECT  15.970 1.980 16.050 2.220 ;
        RECT  15.650 1.820 15.970 2.220 ;
        RECT  13.450 1.820 15.650 2.060 ;
        RECT  14.810 0.750 15.050 1.460 ;
        RECT  14.650 1.060 14.810 1.460 ;
        RECT  12.620 3.080 14.210 3.320 ;
        RECT  13.210 1.320 13.450 2.060 ;
        RECT  11.800 0.670 13.330 0.910 ;
        RECT  12.620 1.820 13.210 2.060 ;
        RECT  12.380 1.820 12.620 3.320 ;
        RECT  12.220 2.250 12.380 2.650 ;
        RECT  11.680 1.460 12.100 1.700 ;
        RECT  11.480 0.670 11.800 1.120 ;
        RECT  11.440 1.460 11.680 3.380 ;
        RECT  11.400 0.860 11.480 1.120 ;
        RECT  10.350 1.460 11.440 1.700 ;
        RECT  11.200 2.980 11.440 3.380 ;
        RECT  9.770 0.860 11.400 1.100 ;
        RECT  10.110 1.460 10.350 2.760 ;
        RECT  9.530 0.860 9.770 3.270 ;
        RECT  9.310 3.550 9.710 3.850 ;
        RECT  9.010 0.890 9.530 1.130 ;
        RECT  8.960 3.030 9.530 3.270 ;
        RECT  8.260 3.550 9.310 3.790 ;
        RECT  9.010 1.410 9.250 2.690 ;
        RECT  8.510 1.410 9.010 1.650 ;
        RECT  8.600 2.450 9.010 2.690 ;
        RECT  7.990 1.930 8.730 2.170 ;
        RECT  8.280 2.450 8.600 3.250 ;
        RECT  8.270 1.250 8.510 1.650 ;
        RECT  8.200 2.900 8.280 3.250 ;
        RECT  7.950 3.520 8.260 3.790 ;
        RECT  7.950 1.130 7.990 2.170 ;
        RECT  7.750 1.130 7.950 3.790 ;
        RECT  6.830 1.130 7.750 1.370 ;
        RECT  7.710 1.930 7.750 3.790 ;
        RECT  6.570 2.930 7.710 3.170 ;
        RECT  7.230 1.770 7.470 2.570 ;
        RECT  5.440 1.770 7.230 2.010 ;
        RECT  6.670 1.130 6.830 1.490 ;
        RECT  6.430 0.670 6.670 1.490 ;
        RECT  5.910 2.290 6.460 2.530 ;
        RECT  6.260 0.670 6.430 0.910 ;
        RECT  5.670 2.290 5.910 3.850 ;
        RECT  3.460 3.610 5.670 3.850 ;
        RECT  5.430 1.480 5.440 2.010 ;
        RECT  5.390 1.280 5.430 2.010 ;
        RECT  5.150 1.270 5.390 3.330 ;
        RECT  5.110 1.270 5.150 1.680 ;
        RECT  3.790 3.090 5.150 3.330 ;
        RECT  5.030 1.280 5.110 1.680 ;
        RECT  4.630 2.000 4.870 2.410 ;
        RECT  3.000 2.000 4.630 2.240 ;
        RECT  3.550 2.520 3.790 3.330 ;
        RECT  3.390 2.520 3.550 2.760 ;
        RECT  3.220 3.610 3.460 4.350 ;
        RECT  1.790 4.110 3.220 4.350 ;
        RECT  2.760 1.390 3.000 3.330 ;
        RECT  2.370 1.390 2.760 1.630 ;
        RECT  2.720 3.090 2.760 3.330 ;
        RECT  2.480 3.090 2.720 3.830 ;
        RECT  2.150 1.870 2.390 2.390 ;
        RECT  2.090 1.870 2.150 2.110 ;
        RECT  1.850 1.310 2.090 2.110 ;
        RECT  0.490 1.310 1.850 1.550 ;
        RECT  1.550 3.260 1.790 4.350 ;
        RECT  0.490 3.260 1.550 3.500 ;
        RECT  0.400 1.310 0.490 1.790 ;
        RECT  0.400 3.100 0.490 3.500 ;
        RECT  0.250 1.310 0.400 3.500 ;
        RECT  0.160 1.320 0.250 3.500 ;
    END
END DFFSRHQX1

MACRO DFFSRXL
    CLASS CORE ;
    FOREIGN DFFSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.510 3.940 4.910 4.370 ;
        RECT  4.910 3.940 5.890 4.180 ;
        RECT  5.890 3.940 6.130 4.360 ;
        RECT  6.130 4.080 6.150 4.360 ;
        RECT  6.150 4.120 7.780 4.360 ;
        RECT  7.780 4.120 8.130 4.370 ;
        RECT  8.130 4.130 11.420 4.370 ;
        RECT  11.420 4.070 11.430 4.370 ;
        RECT  11.430 4.030 11.670 4.370 ;
        RECT  11.670 4.030 11.680 4.330 ;
        RECT  11.680 4.030 12.090 4.270 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.140 1.830 6.150 2.120 ;
        RECT  6.150 1.710 6.490 2.120 ;
        RECT  6.490 1.710 6.610 2.110 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.070 0.680 14.310 4.190 ;
        RECT  14.310 3.950 14.410 4.320 ;
        RECT  14.410 3.950 14.570 4.340 ;
        RECT  14.310 0.680 14.910 0.920 ;
        RECT  14.570 3.950 14.970 4.350 ;
        RECT  14.970 4.070 14.980 4.330 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.040 2.950 16.210 3.210 ;
        RECT  16.210 2.950 16.250 4.350 ;
        RECT  16.250 0.680 16.620 4.350 ;
        RECT  16.620 0.680 16.680 0.920 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.580 2.390 1.590 2.660 ;
        RECT  1.590 2.390 1.990 2.700 ;
        RECT  1.990 2.390 2.440 2.660 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  7.980 2.360 8.580 2.710 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.880 5.440 ;
        RECT  0.880 4.240 0.890 5.440 ;
        RECT  0.890 4.120 1.290 5.440 ;
        RECT  1.290 4.240 1.300 5.440 ;
        RECT  1.300 4.640 3.610 5.440 ;
        RECT  3.610 4.480 4.010 5.440 ;
        RECT  4.010 4.640 5.210 5.440 ;
        RECT  5.210 4.480 5.610 5.440 ;
        RECT  8.530 3.510 8.690 3.750 ;
        RECT  8.690 3.510 8.930 3.850 ;
        RECT  8.930 3.610 10.720 3.850 ;
        RECT  10.720 3.360 10.960 3.850 ;
        RECT  5.610 4.640 12.420 5.440 ;
        RECT  10.960 3.360 12.420 3.600 ;
        RECT  12.420 3.360 12.660 5.440 ;
        RECT  12.660 4.640 13.270 5.440 ;
        RECT  13.270 3.580 13.670 5.440 ;
        RECT  13.670 4.640 15.380 5.440 ;
        RECT  15.380 3.980 15.390 5.440 ;
        RECT  15.390 3.490 15.790 5.440 ;
        RECT  15.790 3.980 15.800 5.440 ;
        RECT  15.800 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  1.090 1.420 1.750 1.660 ;
        RECT  0.000 -0.400 1.750 0.400 ;
        RECT  1.750 -0.400 1.990 1.660 ;
        RECT  1.990 -0.400 3.620 0.400 ;
        RECT  3.620 -0.400 3.630 0.730 ;
        RECT  3.630 -0.400 4.030 0.850 ;
        RECT  4.030 -0.400 4.040 0.730 ;
        RECT  4.040 -0.400 6.830 0.400 ;
        RECT  6.830 -0.400 7.230 0.850 ;
        RECT  7.230 -0.400 8.920 0.400 ;
        RECT  8.920 -0.400 9.320 1.570 ;
        RECT  9.320 -0.400 11.540 0.400 ;
        RECT  11.540 -0.400 11.550 1.290 ;
        RECT  11.550 -0.400 11.950 1.410 ;
        RECT  11.950 -0.400 11.960 1.290 ;
        RECT  11.960 -0.400 15.380 0.400 ;
        RECT  15.380 -0.400 15.390 1.430 ;
        RECT  15.390 -0.400 15.790 1.630 ;
        RECT  15.790 -0.400 15.800 1.430 ;
        RECT  15.800 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.830 1.910 15.940 2.150 ;
        RECT  14.590 1.340 14.830 3.430 ;
        RECT  13.550 1.260 13.790 3.080 ;
        RECT  13.090 1.260 13.550 1.500 ;
        RECT  11.250 2.840 13.550 3.080 ;
        RECT  12.550 2.210 12.710 2.450 ;
        RECT  12.310 1.850 12.550 2.450 ;
        RECT  10.610 1.850 12.310 2.090 ;
        RECT  10.850 2.790 11.250 3.080 ;
        RECT  9.920 0.680 10.930 0.920 ;
        RECT  10.440 1.330 10.610 2.090 ;
        RECT  10.200 1.330 10.440 3.330 ;
        RECT  9.810 3.090 10.200 3.330 ;
        RECT  9.680 0.680 9.920 2.760 ;
        RECT  8.440 1.850 9.680 2.090 ;
        RECT  9.530 2.520 9.680 2.760 ;
        RECT  9.290 2.520 9.530 3.220 ;
        RECT  8.090 2.980 9.290 3.220 ;
        RECT  8.200 1.490 8.440 2.090 ;
        RECT  7.750 0.780 8.240 1.020 ;
        RECT  8.030 1.490 8.200 1.730 ;
        RECT  7.850 2.980 8.090 3.840 ;
        RECT  6.650 3.600 7.850 3.840 ;
        RECT  7.510 0.780 7.750 1.370 ;
        RECT  6.550 1.130 7.510 1.370 ;
        RECT  7.120 2.430 7.330 3.320 ;
        RECT  7.120 1.650 7.280 1.890 ;
        RECT  6.930 1.650 7.120 3.320 ;
        RECT  6.880 1.650 6.930 3.140 ;
        RECT  5.870 2.900 6.880 3.140 ;
        RECT  6.410 3.420 6.650 3.840 ;
        RECT  6.310 0.750 6.550 1.370 ;
        RECT  3.960 3.420 6.410 3.660 ;
        RECT  5.350 0.750 6.310 0.990 ;
        RECT  5.630 2.430 5.870 3.140 ;
        RECT  5.110 0.750 5.350 3.140 ;
        RECT  3.590 2.900 5.110 3.140 ;
        RECT  4.430 2.210 4.830 2.570 ;
        RECT  3.070 2.210 4.430 2.450 ;
        RECT  3.720 3.420 3.960 3.840 ;
        RECT  3.090 3.600 3.720 3.840 ;
        RECT  3.350 2.740 3.590 3.140 ;
        RECT  2.690 3.600 3.090 4.370 ;
        RECT  2.830 1.310 3.070 3.320 ;
        RECT  2.370 1.310 2.830 1.550 ;
        RECT  2.250 3.080 2.830 3.320 ;
        RECT  1.270 3.600 2.690 3.840 ;
        RECT  0.530 0.680 1.290 0.920 ;
        RECT  1.070 2.340 1.270 3.840 ;
        RECT  1.030 2.180 1.070 3.840 ;
        RECT  0.830 2.180 1.030 2.580 ;
        RECT  0.530 4.130 0.600 4.370 ;
        RECT  0.530 3.110 0.570 3.510 ;
        RECT  0.290 0.680 0.530 4.370 ;
        RECT  0.200 4.130 0.290 4.370 ;
    END
END DFFSRXL

MACRO DFFSRX4
    CLASS CORE ;
    FOREIGN DFFSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSRXL ;
    SIZE 23.100 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.120 3.990 4.520 4.360 ;
        RECT  4.520 4.120 8.040 4.360 ;
        RECT  8.040 3.940 8.460 4.360 ;
        RECT  8.460 3.940 12.990 4.180 ;
        RECT  12.990 3.940 13.440 4.350 ;
        RECT  13.440 3.940 13.690 4.340 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.010 2.380 6.480 2.810 ;
        RECT  6.480 2.400 6.550 2.800 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  19.910 1.820 20.070 3.220 ;
        RECT  20.070 1.590 20.080 3.220 ;
        RECT  20.080 1.390 20.350 3.220 ;
        RECT  20.350 1.390 20.480 3.150 ;
        RECT  20.480 1.590 20.490 2.950 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.230 1.820 21.610 3.220 ;
        RECT  21.610 1.590 21.620 3.220 ;
        RECT  21.620 1.390 21.670 3.220 ;
        RECT  21.670 1.390 22.020 3.150 ;
        RECT  22.020 1.590 22.030 2.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.210 2.610 1.520 3.200 ;
        RECT  1.520 2.610 1.610 3.210 ;
        RECT  1.610 2.950 1.780 3.210 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.700 1.890 0.860 2.290 ;
        RECT  0.860 1.830 0.940 2.290 ;
        RECT  0.940 1.830 1.110 2.260 ;
        RECT  1.110 1.830 1.120 2.090 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.980 5.440 ;
        RECT  0.980 4.480 1.380 5.440 ;
        RECT  1.380 4.640 3.450 5.440 ;
        RECT  3.450 4.480 3.850 5.440 ;
        RECT  3.850 4.640 8.950 5.440 ;
        RECT  8.950 4.480 9.350 5.440 ;
        RECT  9.350 4.640 11.510 5.440 ;
        RECT  11.510 4.480 11.910 5.440 ;
        RECT  11.910 4.640 14.630 5.440 ;
        RECT  14.630 3.100 15.030 5.440 ;
        RECT  15.030 4.640 16.600 5.440 ;
        RECT  16.600 3.810 16.610 5.440 ;
        RECT  16.610 3.610 17.010 5.440 ;
        RECT  17.010 3.810 17.020 5.440 ;
        RECT  17.020 4.640 19.460 5.440 ;
        RECT  19.460 4.210 19.470 5.440 ;
        RECT  19.470 4.010 19.870 5.440 ;
        RECT  19.870 4.210 19.880 5.440 ;
        RECT  19.880 4.640 20.870 5.440 ;
        RECT  20.870 4.210 20.880 5.440 ;
        RECT  20.880 4.010 21.280 5.440 ;
        RECT  21.280 4.210 21.290 5.440 ;
        RECT  21.290 4.640 22.280 5.440 ;
        RECT  22.280 4.210 22.290 5.440 ;
        RECT  22.290 4.010 22.690 5.440 ;
        RECT  22.690 4.210 22.700 5.440 ;
        RECT  22.700 4.640 23.100 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.910 0.400 ;
        RECT  0.910 -0.400 1.310 0.560 ;
        RECT  1.310 -0.400 3.220 0.400 ;
        RECT  3.220 -0.400 3.230 0.730 ;
        RECT  3.230 -0.400 3.630 0.850 ;
        RECT  3.630 -0.400 3.640 0.730 ;
        RECT  3.640 -0.400 6.040 0.400 ;
        RECT  6.040 -0.400 6.050 0.800 ;
        RECT  6.050 -0.400 6.450 0.920 ;
        RECT  6.450 -0.400 6.460 0.800 ;
        RECT  6.460 -0.400 8.930 0.400 ;
        RECT  8.930 -0.400 9.170 1.400 ;
        RECT  9.170 -0.400 11.340 0.400 ;
        RECT  11.340 -0.400 11.350 0.820 ;
        RECT  11.350 -0.400 11.750 0.940 ;
        RECT  11.750 -0.400 11.760 0.820 ;
        RECT  11.760 -0.400 14.280 0.400 ;
        RECT  14.280 -0.400 14.290 0.880 ;
        RECT  14.290 -0.400 14.690 1.080 ;
        RECT  14.690 -0.400 14.700 0.880 ;
        RECT  14.700 -0.400 19.460 0.400 ;
        RECT  19.460 -0.400 19.470 0.910 ;
        RECT  19.470 -0.400 19.870 1.110 ;
        RECT  19.870 -0.400 19.880 0.910 ;
        RECT  19.880 -0.400 20.870 0.400 ;
        RECT  20.870 -0.400 20.880 0.950 ;
        RECT  20.880 -0.400 21.280 1.150 ;
        RECT  21.280 -0.400 21.290 0.950 ;
        RECT  21.290 -0.400 22.280 0.400 ;
        RECT  22.280 -0.400 22.290 0.910 ;
        RECT  22.290 -0.400 22.690 1.110 ;
        RECT  22.690 -0.400 22.700 0.910 ;
        RECT  22.700 -0.400 23.100 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  22.360 2.170 22.600 3.730 ;
        RECT  19.640 3.490 22.360 3.730 ;
        RECT  19.400 1.550 19.640 3.730 ;
        RECT  18.930 1.550 19.400 1.790 ;
        RECT  18.610 3.330 19.400 3.730 ;
        RECT  18.720 2.130 19.120 2.530 ;
        RECT  18.690 1.390 18.930 1.790 ;
        RECT  18.410 2.140 18.720 2.530 ;
        RECT  18.090 0.680 18.490 0.960 ;
        RECT  18.210 1.480 18.410 3.050 ;
        RECT  18.170 1.480 18.210 3.640 ;
        RECT  17.730 1.480 18.170 1.720 ;
        RECT  17.970 2.810 18.170 3.640 ;
        RECT  16.970 0.680 18.090 0.920 ;
        RECT  17.810 3.080 17.970 3.640 ;
        RECT  17.650 2.060 17.890 2.460 ;
        RECT  15.790 3.080 17.810 3.320 ;
        RECT  17.330 1.200 17.730 1.720 ;
        RECT  13.300 2.060 17.650 2.300 ;
        RECT  16.210 1.480 17.330 1.720 ;
        RECT  16.730 0.680 16.970 1.200 ;
        RECT  16.570 0.720 16.730 1.200 ;
        RECT  15.450 0.720 16.570 0.960 ;
        RECT  15.810 1.240 16.210 1.720 ;
        RECT  15.630 3.080 15.790 3.630 ;
        RECT  15.390 2.580 15.630 3.630 ;
        RECT  15.290 0.720 15.450 1.320 ;
        RECT  14.270 2.580 15.390 2.820 ;
        RECT  15.210 0.720 15.290 1.610 ;
        RECT  15.050 0.920 15.210 1.610 ;
        RECT  13.850 1.370 15.050 1.610 ;
        RECT  14.110 3.420 14.350 4.370 ;
        RECT  14.030 2.580 14.270 3.140 ;
        RECT  7.860 3.420 14.110 3.660 ;
        RECT  13.870 2.860 14.030 3.140 ;
        RECT  12.180 2.900 13.870 3.140 ;
        RECT  13.610 0.940 13.850 1.610 ;
        RECT  13.060 0.830 13.300 2.300 ;
        RECT  12.690 0.830 13.060 1.070 ;
        RECT  12.870 1.920 13.060 2.300 ;
        RECT  12.460 1.920 12.870 2.620 ;
        RECT  11.630 1.400 12.770 1.640 ;
        RECT  10.910 1.920 12.460 2.160 ;
        RECT  11.940 2.440 12.180 3.140 ;
        RECT  11.780 2.440 11.940 2.680 ;
        RECT  11.390 1.220 11.630 1.640 ;
        RECT  10.930 1.220 11.390 1.460 ;
        RECT  10.690 0.670 10.930 1.460 ;
        RECT  10.670 1.750 10.910 3.140 ;
        RECT  9.870 0.670 10.690 0.910 ;
        RECT  10.390 1.750 10.670 1.990 ;
        RECT  10.230 2.900 10.670 3.140 ;
        RECT  10.150 1.190 10.390 1.990 ;
        RECT  9.870 2.270 10.390 2.510 ;
        RECT  9.630 0.670 9.870 2.510 ;
        RECT  9.060 2.270 9.630 2.510 ;
        RECT  8.820 2.040 9.060 2.510 ;
        RECT  8.650 2.040 8.820 2.280 ;
        RECT  8.380 2.900 8.540 3.140 ;
        RECT  8.350 2.560 8.380 3.140 ;
        RECT  8.140 1.370 8.350 3.140 ;
        RECT  7.100 0.770 8.230 1.010 ;
        RECT  8.110 1.370 8.140 2.800 ;
        RECT  7.510 2.020 8.110 2.260 ;
        RECT  7.620 3.080 7.860 3.660 ;
        RECT  7.150 3.080 7.620 3.320 ;
        RECT  5.040 3.600 7.340 3.840 ;
        RECT  6.910 1.720 7.150 3.320 ;
        RECT  6.860 0.770 7.100 1.440 ;
        RECT  6.750 1.720 6.910 1.960 ;
        RECT  5.730 3.080 6.910 3.320 ;
        RECT  5.210 1.200 6.860 1.440 ;
        RECT  5.490 2.370 5.730 3.320 ;
        RECT  4.970 1.200 5.210 3.100 ;
        RECT  4.800 3.470 5.040 3.840 ;
        RECT  4.710 1.200 4.970 1.440 ;
        RECT  4.790 2.860 4.970 3.100 ;
        RECT  3.160 3.470 4.800 3.710 ;
        RECT  4.390 2.860 4.790 3.190 ;
        RECT  4.490 1.870 4.730 2.270 ;
        RECT  4.420 1.870 4.490 2.110 ;
        RECT  4.180 1.690 4.420 2.110 ;
        RECT  3.410 2.860 4.390 3.100 ;
        RECT  2.880 1.690 4.180 1.930 ;
        RECT  3.170 2.210 3.410 3.100 ;
        RECT  2.920 3.470 3.160 4.100 ;
        RECT  0.570 3.860 2.920 4.100 ;
        RECT  2.640 1.190 2.880 2.660 ;
        RECT  2.110 1.190 2.640 1.430 ;
        RECT  2.490 2.420 2.640 2.660 ;
        RECT  2.250 2.420 2.490 3.570 ;
        RECT  1.950 1.710 2.190 2.140 ;
        RECT  1.770 1.710 1.950 1.950 ;
        RECT  1.530 1.310 1.770 1.950 ;
        RECT  0.570 1.310 1.530 1.550 ;
        RECT  0.460 1.150 0.570 1.550 ;
        RECT  0.460 3.440 0.570 4.100 ;
        RECT  0.330 1.150 0.460 4.100 ;
        RECT  0.220 1.150 0.330 3.840 ;
        RECT  0.170 1.150 0.220 1.550 ;
        RECT  0.170 3.440 0.220 3.840 ;
    END
END DFFSRX4

MACRO DFFSRX2
    CLASS CORE ;
    FOREIGN DFFSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSRXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.070 3.940 4.470 4.370 ;
        RECT  4.470 3.940 5.430 4.180 ;
        RECT  5.430 3.940 5.670 4.360 ;
        RECT  5.670 4.120 7.570 4.360 ;
        RECT  7.570 4.120 7.810 4.370 ;
        RECT  7.810 4.130 11.010 4.370 ;
        RECT  11.010 4.080 11.160 4.370 ;
        RECT  11.160 4.030 11.560 4.370 ;
        RECT  11.560 4.030 11.670 4.330 ;
        RECT  11.670 4.070 11.680 4.330 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.480 1.770 5.490 2.090 ;
        RECT  5.490 1.770 5.880 2.100 ;
        RECT  5.880 1.770 5.980 2.180 ;
        RECT  5.980 1.780 6.120 2.180 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.530 2.890 14.630 3.290 ;
        RECT  14.630 2.660 14.730 3.290 ;
        RECT  14.730 2.640 14.780 3.290 ;
        RECT  14.780 1.150 14.930 3.290 ;
        RECT  14.930 1.150 14.980 3.210 ;
        RECT  14.980 1.150 15.020 3.130 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.380 1.260 15.970 1.540 ;
        RECT  15.930 2.890 16.090 3.290 ;
        RECT  15.970 1.150 16.090 1.550 ;
        RECT  16.090 1.150 16.330 3.290 ;
        RECT  16.330 1.150 16.370 1.550 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.340 2.380 1.870 2.820 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  7.460 2.250 8.210 2.720 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.020 5.440 ;
        RECT  1.020 4.480 1.420 5.440 ;
        RECT  1.420 4.640 3.390 5.440 ;
        RECT  3.390 4.480 3.790 5.440 ;
        RECT  3.790 4.640 4.750 5.440 ;
        RECT  4.750 4.480 5.150 5.440 ;
        RECT  8.250 3.510 8.650 3.850 ;
        RECT  8.650 3.610 10.460 3.850 ;
        RECT  10.460 3.460 10.700 3.850 ;
        RECT  5.150 4.640 12.070 5.440 ;
        RECT  10.700 3.460 12.070 3.700 ;
        RECT  12.070 3.460 12.310 5.440 ;
        RECT  12.310 4.640 13.010 5.440 ;
        RECT  13.010 3.730 13.020 5.440 ;
        RECT  13.020 3.530 13.420 5.440 ;
        RECT  13.420 3.730 13.430 5.440 ;
        RECT  13.430 4.640 15.310 5.440 ;
        RECT  15.310 4.350 15.320 5.440 ;
        RECT  15.320 4.150 15.720 5.440 ;
        RECT  15.720 4.350 15.730 5.440 ;
        RECT  15.730 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.440 0.400 ;
        RECT  0.440 -0.400 0.840 0.560 ;
        RECT  0.840 -0.400 3.230 0.400 ;
        RECT  3.230 -0.400 3.240 0.890 ;
        RECT  3.240 -0.400 3.640 1.090 ;
        RECT  3.640 -0.400 3.650 0.890 ;
        RECT  3.650 -0.400 6.310 0.400 ;
        RECT  6.310 -0.400 6.710 0.910 ;
        RECT  6.710 -0.400 8.340 0.400 ;
        RECT  8.340 -0.400 8.350 1.210 ;
        RECT  8.350 -0.400 8.750 1.410 ;
        RECT  8.750 -0.400 8.760 1.210 ;
        RECT  8.760 -0.400 10.870 0.400 ;
        RECT  10.870 -0.400 11.270 0.560 ;
        RECT  11.270 -0.400 13.930 0.400 ;
        RECT  13.930 -0.400 14.330 0.560 ;
        RECT  14.330 -0.400 15.340 0.400 ;
        RECT  15.340 -0.400 15.350 0.670 ;
        RECT  15.350 -0.400 15.750 0.870 ;
        RECT  15.750 -0.400 15.760 0.670 ;
        RECT  15.760 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  15.650 2.180 15.810 2.580 ;
        RECT  15.410 2.180 15.650 3.870 ;
        RECT  14.270 3.630 15.410 3.870 ;
        RECT  14.250 1.530 14.320 1.930 ;
        RECT  14.250 3.630 14.270 4.120 ;
        RECT  14.010 1.530 14.250 4.120 ;
        RECT  13.920 1.530 14.010 1.930 ;
        RECT  13.870 3.720 14.010 4.120 ;
        RECT  13.640 2.210 13.730 2.610 ;
        RECT  13.400 1.270 13.640 3.170 ;
        RECT  13.520 0.730 13.600 0.970 ;
        RECT  13.200 0.730 13.520 0.980 ;
        RECT  12.440 1.270 13.400 1.510 ;
        RECT  10.960 2.930 13.400 3.170 ;
        RECT  12.080 0.740 13.200 0.980 ;
        RECT  12.090 1.850 12.330 2.260 ;
        RECT  10.210 1.850 12.090 2.090 ;
        RECT  11.760 0.740 12.080 1.150 ;
        RECT  11.680 0.750 11.760 1.150 ;
        RECT  10.720 2.370 10.960 3.170 ;
        RECT  10.560 2.370 10.720 2.610 ;
        RECT  9.270 0.730 10.460 0.970 ;
        RECT  10.170 1.330 10.210 2.090 ;
        RECT  9.930 1.330 10.170 3.330 ;
        RECT  9.630 1.330 9.930 1.570 ;
        RECT  9.550 3.090 9.930 3.330 ;
        RECT  9.270 2.520 9.650 2.760 ;
        RECT  9.030 0.730 9.270 3.230 ;
        RECT  7.870 1.690 9.030 1.930 ;
        RECT  7.890 2.990 9.030 3.230 ;
        RECT  7.650 2.990 7.890 3.840 ;
        RECT  7.470 1.360 7.870 1.930 ;
        RECT  7.190 0.770 7.730 1.010 ;
        RECT  7.490 3.440 7.650 3.840 ;
        RECT  6.190 3.600 7.490 3.840 ;
        RECT  6.950 0.770 7.190 1.390 ;
        RECT  6.860 1.650 7.100 3.320 ;
        RECT  5.100 1.150 6.950 1.390 ;
        RECT  6.400 1.650 6.860 1.890 ;
        RECT  6.470 2.900 6.860 3.320 ;
        RECT  5.620 2.900 6.470 3.140 ;
        RECT  5.950 3.420 6.190 3.840 ;
        RECT  2.860 3.420 5.950 3.660 ;
        RECT  5.380 2.510 5.620 3.140 ;
        RECT  4.860 1.150 5.100 3.020 ;
        RECT  4.780 1.150 4.860 1.390 ;
        RECT  3.620 2.780 4.860 3.020 ;
        RECT  4.340 1.660 4.580 2.060 ;
        RECT  2.600 1.820 4.340 2.060 ;
        RECT  3.220 2.780 3.620 3.140 ;
        RECT  2.860 4.130 2.940 4.370 ;
        RECT  2.540 3.420 2.860 4.370 ;
        RECT  2.440 1.820 2.600 3.140 ;
        RECT  1.070 3.420 2.540 3.660 ;
        RECT  2.200 0.750 2.440 3.140 ;
        RECT  2.160 4.130 2.220 4.370 ;
        RECT  1.820 3.940 2.160 4.370 ;
        RECT  1.300 0.690 1.920 0.930 ;
        RECT  0.490 3.940 1.820 4.180 ;
        RECT  1.060 0.690 1.300 1.630 ;
        RECT  0.830 2.670 1.070 3.660 ;
        RECT  0.570 1.390 1.060 1.630 ;
        RECT  0.740 2.670 0.830 3.070 ;
        RECT  0.410 1.390 0.570 1.790 ;
        RECT  0.410 3.350 0.490 4.180 ;
        RECT  0.250 1.390 0.410 4.180 ;
        RECT  0.170 1.390 0.250 3.590 ;
    END
END DFFSRX2

MACRO DFFSRX1
    CLASS CORE ;
    FOREIGN DFFSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSRXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.590 3.940 4.990 4.350 ;
        RECT  4.990 3.940 5.970 4.180 ;
        RECT  5.970 3.940 6.210 4.360 ;
        RECT  6.210 4.120 8.130 4.360 ;
        RECT  8.130 4.120 8.370 4.370 ;
        RECT  8.370 4.130 11.670 4.370 ;
        RECT  11.670 4.080 11.720 4.370 ;
        RECT  11.720 4.030 11.960 4.370 ;
        RECT  11.960 4.030 12.080 4.340 ;
        RECT  12.080 4.030 12.120 4.330 ;
        RECT  12.120 4.070 12.340 4.330 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.130 1.820 6.540 2.190 ;
        RECT  6.540 1.780 6.780 2.190 ;
        RECT  6.780 1.820 6.790 2.190 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.410 0.730 14.650 3.750 ;
        RECT  14.650 3.510 14.720 3.750 ;
        RECT  14.720 3.510 14.910 3.770 ;
        RECT  14.910 3.510 14.980 4.150 ;
        RECT  14.980 3.530 15.150 4.150 ;
        RECT  15.150 3.750 15.310 4.150 ;
        RECT  14.650 0.730 15.310 0.970 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.040 2.950 16.150 3.210 ;
        RECT  16.150 2.950 16.560 3.220 ;
        RECT  16.560 2.950 16.720 3.430 ;
        RECT  16.570 1.190 16.720 1.590 ;
        RECT  16.720 1.190 16.960 3.430 ;
        RECT  16.960 1.190 16.970 1.590 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 2.380 1.930 2.830 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  8.120 2.330 8.760 2.720 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.190 5.440 ;
        RECT  1.190 4.480 1.590 5.440 ;
        RECT  1.590 4.640 3.910 5.440 ;
        RECT  3.910 4.480 4.310 5.440 ;
        RECT  4.310 4.640 5.290 5.440 ;
        RECT  5.290 4.480 5.690 5.440 ;
        RECT  8.810 3.510 8.970 3.750 ;
        RECT  8.970 3.510 9.210 3.850 ;
        RECT  9.210 3.610 11.010 3.850 ;
        RECT  11.010 3.460 11.250 3.850 ;
        RECT  5.690 4.640 12.700 5.440 ;
        RECT  11.250 3.460 12.700 3.700 ;
        RECT  12.700 3.460 12.940 5.440 ;
        RECT  12.940 4.640 13.540 5.440 ;
        RECT  13.540 3.580 13.550 5.440 ;
        RECT  13.550 3.460 13.950 5.440 ;
        RECT  13.950 3.580 13.960 5.440 ;
        RECT  13.960 4.640 15.720 5.440 ;
        RECT  15.720 3.460 16.120 5.440 ;
        RECT  16.120 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.170 0.400 ;
        RECT  1.170 -0.400 1.180 1.330 ;
        RECT  1.180 -0.400 1.580 1.450 ;
        RECT  1.580 -0.400 1.590 1.330 ;
        RECT  1.590 -0.400 3.890 0.400 ;
        RECT  3.890 -0.400 3.900 0.730 ;
        RECT  3.900 -0.400 4.300 0.930 ;
        RECT  4.300 -0.400 4.310 0.730 ;
        RECT  4.310 -0.400 6.840 0.400 ;
        RECT  6.840 -0.400 7.240 0.850 ;
        RECT  7.240 -0.400 8.930 0.400 ;
        RECT  8.930 -0.400 9.330 1.540 ;
        RECT  9.330 -0.400 11.480 0.400 ;
        RECT  11.480 -0.400 11.880 0.560 ;
        RECT  11.880 -0.400 15.720 0.400 ;
        RECT  15.720 -0.400 15.730 0.990 ;
        RECT  15.730 -0.400 16.130 1.480 ;
        RECT  16.130 -0.400 16.140 0.990 ;
        RECT  16.140 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.080 1.870 16.480 2.270 ;
        RECT  15.170 1.950 16.080 2.190 ;
        RECT  14.930 1.390 15.170 3.170 ;
        RECT  13.890 0.780 14.130 1.510 ;
        RECT  13.450 2.250 14.070 2.650 ;
        RECT  12.690 0.780 13.890 1.020 ;
        RECT  13.210 1.310 13.450 3.170 ;
        RECT  13.050 1.310 13.210 1.550 ;
        RECT  11.550 2.930 13.210 3.170 ;
        RECT  12.650 1.850 12.890 2.260 ;
        RECT  12.450 0.780 12.690 1.510 ;
        RECT  10.770 1.850 12.650 2.090 ;
        RECT  12.290 1.110 12.450 1.510 ;
        RECT  11.310 2.680 11.550 3.170 ;
        RECT  11.140 2.680 11.310 2.920 ;
        RECT  9.920 0.730 11.050 0.970 ;
        RECT  10.730 1.300 10.770 2.090 ;
        RECT  10.490 1.300 10.730 3.330 ;
        RECT  10.200 1.300 10.490 1.540 ;
        RECT  10.110 3.090 10.490 3.330 ;
        RECT  9.910 2.520 10.210 2.760 ;
        RECT  9.910 0.730 9.920 2.060 ;
        RECT  9.830 0.730 9.910 2.760 ;
        RECT  9.670 0.730 9.830 3.230 ;
        RECT  9.590 1.820 9.670 3.230 ;
        RECT  9.580 1.820 9.590 2.590 ;
        RECT  8.450 2.990 9.590 3.230 ;
        RECT  8.450 1.820 9.580 2.060 ;
        RECT  8.210 1.460 8.450 2.060 ;
        RECT  8.370 2.990 8.450 3.830 ;
        RECT  8.210 2.990 8.370 3.840 ;
        RECT  7.770 0.770 8.280 1.010 ;
        RECT  8.050 1.460 8.210 1.700 ;
        RECT  8.050 3.430 8.210 3.840 ;
        RECT  6.730 3.600 8.050 3.840 ;
        RECT  7.530 0.770 7.770 1.370 ;
        RECT  5.840 1.130 7.530 1.370 ;
        RECT  7.460 2.430 7.500 3.320 ;
        RECT  7.220 1.650 7.460 3.320 ;
        RECT  7.050 1.650 7.220 1.890 ;
        RECT  7.010 2.900 7.220 3.320 ;
        RECT  6.280 2.900 7.010 3.140 ;
        RECT  6.490 3.420 6.730 3.840 ;
        RECT  4.260 3.420 6.490 3.660 ;
        RECT  6.040 2.510 6.280 3.140 ;
        RECT  5.760 1.090 5.840 1.490 ;
        RECT  5.520 1.090 5.760 3.140 ;
        RECT  5.440 1.090 5.520 1.490 ;
        RECT  4.080 2.900 5.520 3.140 ;
        RECT  5.000 1.780 5.240 2.180 ;
        RECT  3.500 1.940 5.000 2.180 ;
        RECT  4.020 3.420 4.260 4.120 ;
        RECT  3.840 2.460 4.080 3.140 ;
        RECT  3.310 3.880 4.020 4.120 ;
        RECT  3.260 1.220 3.500 3.100 ;
        RECT  3.070 3.420 3.310 4.120 ;
        RECT  2.920 1.220 3.260 1.460 ;
        RECT  2.740 2.860 3.260 3.100 ;
        RECT  1.100 3.420 3.070 3.660 ;
        RECT  2.740 1.740 2.980 2.140 ;
        RECT  2.520 1.060 2.920 1.460 ;
        RECT  0.700 1.740 2.740 1.980 ;
        RECT  0.580 3.940 2.630 4.180 ;
        RECT  0.860 2.450 1.100 3.660 ;
        RECT  0.580 1.320 0.700 1.980 ;
        RECT  0.340 1.320 0.580 4.180 ;
        RECT  0.300 1.320 0.340 1.720 ;
    END
END DFFSRX1

MACRO DFFSHQXL
    CLASS CORE ;
    FOREIGN DFFSHQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.290 2.530 4.820 2.930 ;
        RECT  4.820 2.390 5.080 2.930 ;
        RECT  5.080 2.650 5.170 2.930 ;
        RECT  5.170 2.690 5.300 2.930 ;
        RECT  5.300 2.690 5.540 4.180 ;
        RECT  5.540 3.940 7.160 4.180 ;
        RECT  7.160 3.940 7.400 4.370 ;
        RECT  7.400 4.080 7.470 4.370 ;
        RECT  7.470 4.130 11.010 4.370 ;
        RECT  11.010 4.080 11.150 4.370 ;
        RECT  11.150 2.240 11.290 4.370 ;
        RECT  11.290 2.080 11.390 4.370 ;
        RECT  11.390 2.080 11.430 2.640 ;
        RECT  11.430 2.080 11.690 2.480 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.830 3.220 11.990 3.620 ;
        RECT  11.990 2.790 12.230 3.620 ;
        RECT  12.230 2.790 12.650 3.030 ;
        RECT  12.650 2.660 12.750 3.030 ;
        RECT  12.740 1.830 12.750 2.090 ;
        RECT  12.710 1.000 12.750 1.400 ;
        RECT  12.750 1.000 12.990 3.030 ;
        RECT  12.990 1.830 13.000 2.090 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.300 1.270 1.780 1.950 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.770 2.390 1.340 2.890 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.210 5.440 ;
        RECT  1.210 4.480 1.610 5.440 ;
        RECT  1.610 4.640 4.050 5.440 ;
        RECT  4.050 4.090 5.030 5.440 ;
        RECT  5.030 4.640 6.470 5.440 ;
        RECT  6.470 4.480 6.870 5.440 ;
        RECT  6.870 4.640 11.670 5.440 ;
        RECT  11.670 4.480 12.070 5.440 ;
        RECT  12.070 4.640 12.580 5.440 ;
        RECT  12.580 3.510 12.590 5.440 ;
        RECT  12.590 3.310 12.990 5.440 ;
        RECT  12.990 3.510 13.000 5.440 ;
        RECT  13.000 4.640 13.200 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.090 0.400 ;
        RECT  1.090 -0.400 1.490 0.870 ;
        RECT  1.490 -0.400 3.700 0.400 ;
        RECT  3.700 -0.400 3.710 0.730 ;
        RECT  3.710 -0.400 4.110 0.850 ;
        RECT  4.110 -0.400 4.120 0.730 ;
        RECT  4.120 -0.400 6.750 0.400 ;
        RECT  6.750 -0.400 6.990 1.300 ;
        RECT  6.990 -0.400 9.710 0.400 ;
        RECT  9.710 -0.400 10.110 0.560 ;
        RECT  10.110 -0.400 11.350 0.400 ;
        RECT  11.350 -0.400 11.750 0.560 ;
        RECT  11.750 -0.400 13.200 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.130 1.280 12.370 2.510 ;
        RECT  11.130 1.280 12.130 1.520 ;
        RECT  10.890 0.860 11.130 1.520 ;
        RECT  10.790 0.860 10.890 1.100 ;
        RECT  9.970 3.590 10.810 3.830 ;
        RECT  10.390 0.690 10.790 1.100 ;
        RECT  9.870 0.860 10.390 1.100 ;
        RECT  10.150 1.380 10.390 2.710 ;
        RECT  9.970 2.470 10.150 2.710 ;
        RECT  9.730 2.470 9.970 3.830 ;
        RECT  9.630 0.860 9.870 2.190 ;
        RECT  9.430 0.860 9.630 1.100 ;
        RECT  9.450 1.950 9.630 2.190 ;
        RECT  9.210 1.950 9.450 3.130 ;
        RECT  9.140 0.780 9.430 1.100 ;
        RECT  8.220 2.890 9.210 3.130 ;
        RECT  6.810 3.410 9.190 3.650 ;
        RECT  8.370 0.780 9.140 1.020 ;
        RECT  8.800 1.380 9.090 1.620 ;
        RECT  8.560 1.380 8.800 2.370 ;
        RECT  7.850 2.130 8.560 2.370 ;
        RECT  7.790 1.010 7.950 1.410 ;
        RECT  7.610 2.130 7.850 2.610 ;
        RECT  7.550 1.010 7.790 1.840 ;
        RECT  7.330 2.890 7.740 3.130 ;
        RECT  7.330 1.600 7.550 1.840 ;
        RECT  7.090 1.600 7.330 3.130 ;
        RECT  6.570 1.580 6.810 3.650 ;
        RECT  6.470 1.580 6.570 1.820 ;
        RECT  5.870 3.410 6.570 3.650 ;
        RECT  6.230 1.360 6.470 1.820 ;
        RECT  6.090 2.110 6.330 2.690 ;
        RECT  6.110 1.360 6.230 1.600 ;
        RECT  5.870 0.670 6.110 1.600 ;
        RECT  5.950 2.110 6.090 2.350 ;
        RECT  5.710 1.870 5.950 2.350 ;
        RECT  5.470 0.670 5.870 0.910 ;
        RECT  5.450 1.870 5.710 2.110 ;
        RECT  5.210 1.350 5.450 2.110 ;
        RECT  5.050 1.350 5.210 2.080 ;
        RECT  4.770 0.770 5.150 1.010 ;
        RECT  4.050 1.840 5.050 2.080 ;
        RECT  4.050 3.370 4.830 3.610 ;
        RECT  4.530 0.770 4.770 1.370 ;
        RECT  3.290 1.130 4.530 1.370 ;
        RECT  3.810 1.840 4.050 3.610 ;
        RECT  3.530 1.840 3.810 2.080 ;
        RECT  3.290 2.360 3.530 4.050 ;
        RECT  3.250 0.940 3.290 1.370 ;
        RECT  3.250 2.360 3.290 2.600 ;
        RECT  2.550 3.810 3.290 4.050 ;
        RECT  3.010 0.940 3.250 2.600 ;
        RECT  2.370 0.940 3.010 1.180 ;
        RECT  2.780 3.040 3.010 3.440 ;
        RECT  2.450 3.040 2.780 3.450 ;
        RECT  2.400 1.540 2.450 3.450 ;
        RECT  2.210 1.540 2.400 3.440 ;
        RECT  0.790 3.200 2.210 3.440 ;
        RECT  0.490 3.200 0.790 4.020 ;
        RECT  0.490 0.960 0.610 1.360 ;
        RECT  0.390 0.960 0.490 4.020 ;
        RECT  0.250 0.960 0.390 3.440 ;
        RECT  0.210 0.960 0.250 1.360 ;
    END
END DFFSHQXL

MACRO DFFSHQX4
    CLASS CORE ;
    FOREIGN DFFSHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSHQXL ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.490 2.400 4.820 2.880 ;
        RECT  4.820 2.390 5.080 2.880 ;
        RECT  5.080 2.640 5.590 2.880 ;
        RECT  5.590 2.640 5.830 3.660 ;
        RECT  5.830 3.420 7.850 3.660 ;
        RECT  7.850 3.420 8.090 3.730 ;
        RECT  8.090 3.490 9.510 3.730 ;
        RECT  9.510 3.490 9.790 4.180 ;
        RECT  9.790 3.940 14.440 4.180 ;
        RECT  14.440 3.640 14.940 4.180 ;
        RECT  14.940 2.260 14.970 4.180 ;
        RECT  14.970 2.250 15.180 4.180 ;
        RECT  15.180 2.250 15.370 2.660 ;
        RECT  15.370 2.380 16.570 2.660 ;
        RECT  16.570 2.250 16.910 2.660 ;
        RECT  16.910 2.250 16.970 2.650 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.470 0.800 15.870 1.390 ;
        RECT  15.530 3.050 15.930 4.030 ;
        RECT  15.930 3.050 16.170 3.300 ;
        RECT  16.170 3.060 16.930 3.300 ;
        RECT  16.930 2.940 17.050 3.300 ;
        RECT  17.050 2.940 17.270 4.050 ;
        RECT  17.270 2.940 17.710 4.340 ;
        RECT  15.870 1.150 17.910 1.390 ;
        RECT  17.710 2.940 18.070 3.290 ;
        RECT  17.910 0.770 18.070 1.390 ;
        RECT  18.070 0.770 18.310 3.290 ;
        RECT  18.310 3.000 18.320 3.290 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 1.260 1.870 1.730 ;
        RECT  1.870 1.330 1.880 1.730 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.120 1.390 2.660 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.540 5.440 ;
        RECT  1.540 3.900 1.940 5.440 ;
        RECT  1.940 4.640 4.080 5.440 ;
        RECT  4.080 4.480 4.480 5.440 ;
        RECT  4.480 4.640 5.720 5.440 ;
        RECT  5.720 4.480 6.120 5.440 ;
        RECT  6.120 4.640 7.150 5.440 ;
        RECT  7.150 4.060 7.160 5.440 ;
        RECT  7.160 3.940 7.560 5.440 ;
        RECT  7.560 4.060 7.570 5.440 ;
        RECT  7.570 4.640 8.800 5.440 ;
        RECT  8.800 4.130 8.810 5.440 ;
        RECT  8.810 4.010 9.210 5.440 ;
        RECT  9.210 4.130 9.220 5.440 ;
        RECT  9.220 4.640 13.250 5.440 ;
        RECT  13.250 4.480 13.650 5.440 ;
        RECT  13.650 4.640 14.710 5.440 ;
        RECT  14.710 4.480 15.110 5.440 ;
        RECT  15.110 4.640 16.280 5.440 ;
        RECT  16.280 4.090 16.290 5.440 ;
        RECT  16.290 3.600 16.690 5.440 ;
        RECT  16.690 4.090 16.700 5.440 ;
        RECT  16.700 4.640 17.980 5.440 ;
        RECT  17.980 3.600 18.220 5.440 ;
        RECT  18.220 4.640 18.480 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.180 0.400 ;
        RECT  1.180 -0.400 1.190 0.750 ;
        RECT  1.190 -0.400 1.590 0.870 ;
        RECT  1.590 -0.400 1.600 0.750 ;
        RECT  1.600 -0.400 3.780 0.400 ;
        RECT  3.780 -0.400 3.790 0.730 ;
        RECT  3.790 -0.400 4.190 0.850 ;
        RECT  4.190 -0.400 4.200 0.730 ;
        RECT  4.200 -0.400 7.260 0.400 ;
        RECT  7.260 -0.400 7.270 1.320 ;
        RECT  7.270 -0.400 7.670 1.440 ;
        RECT  7.670 -0.400 7.680 1.320 ;
        RECT  7.680 -0.400 8.780 0.400 ;
        RECT  8.780 -0.400 8.790 1.110 ;
        RECT  8.790 -0.400 9.190 1.230 ;
        RECT  9.190 -0.400 9.200 1.110 ;
        RECT  9.200 -0.400 13.020 0.400 ;
        RECT  13.020 -0.400 13.420 0.560 ;
        RECT  13.420 -0.400 14.190 0.400 ;
        RECT  14.190 -0.400 14.590 0.560 ;
        RECT  14.590 -0.400 16.690 0.400 ;
        RECT  16.690 -0.400 17.090 0.870 ;
        RECT  17.090 -0.400 18.480 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  17.630 2.070 17.790 2.470 ;
        RECT  17.390 1.730 17.630 2.470 ;
        RECT  15.020 1.730 17.390 1.970 ;
        RECT  14.780 0.860 15.020 1.970 ;
        RECT  12.240 0.860 14.780 1.100 ;
        RECT  14.210 1.540 14.450 3.290 ;
        RECT  13.540 1.540 14.210 1.780 ;
        RECT  14.050 2.890 14.210 3.290 ;
        RECT  13.710 2.220 13.870 2.620 ;
        RECT  13.470 2.220 13.710 3.660 ;
        RECT  13.120 1.340 13.540 1.780 ;
        RECT  12.230 3.420 13.470 3.660 ;
        RECT  12.720 1.340 13.120 2.350 ;
        RECT  12.230 0.860 12.240 1.630 ;
        RECT  12.080 0.860 12.230 3.660 ;
        RECT  11.990 0.670 12.080 3.660 ;
        RECT  11.840 0.670 11.990 1.630 ;
        RECT  10.390 3.420 11.990 3.660 ;
        RECT  10.720 0.670 11.840 0.910 ;
        RECT  10.750 2.900 11.550 3.140 ;
        RECT  11.320 1.250 11.480 1.490 ;
        RECT  11.080 1.250 11.320 1.750 ;
        RECT  10.750 1.510 11.080 1.750 ;
        RECT  10.510 1.510 10.750 3.140 ;
        RECT  10.480 0.670 10.720 1.230 ;
        RECT  9.960 1.510 10.510 1.750 ;
        RECT  10.030 2.900 10.510 3.140 ;
        RECT  10.320 0.990 10.480 1.230 ;
        RECT  7.670 2.030 10.230 2.270 ;
        RECT  9.630 2.900 10.030 3.210 ;
        RECT  9.950 1.410 9.960 1.750 ;
        RECT  9.550 1.070 9.950 1.750 ;
        RECT  7.990 2.900 9.630 3.140 ;
        RECT  8.430 1.510 9.550 1.750 ;
        RECT  8.110 1.070 8.430 1.750 ;
        RECT  8.030 1.070 8.110 1.470 ;
        RECT  7.430 1.800 7.670 3.140 ;
        RECT  6.940 1.800 7.430 2.040 ;
        RECT  6.600 2.900 7.430 3.140 ;
        RECT  6.350 2.320 7.150 2.560 ;
        RECT  6.830 1.310 6.940 2.040 ;
        RECT  6.700 0.670 6.830 2.040 ;
        RECT  6.400 3.940 6.800 4.370 ;
        RECT  6.590 0.670 6.700 1.630 ;
        RECT  6.180 0.670 6.590 0.910 ;
        RECT  2.490 3.940 6.400 4.180 ;
        RECT  6.110 1.920 6.350 2.560 ;
        RECT  5.680 1.920 6.110 2.160 ;
        RECT  4.790 0.770 5.860 1.010 ;
        RECT  5.530 1.650 5.680 2.160 ;
        RECT  5.440 1.460 5.530 2.160 ;
        RECT  5.130 1.460 5.440 1.890 ;
        RECT  4.200 3.190 5.300 3.430 ;
        RECT  4.200 1.650 5.130 1.890 ;
        RECT  4.550 0.770 4.790 1.370 ;
        RECT  3.270 1.130 4.550 1.370 ;
        RECT  3.960 1.650 4.200 3.430 ;
        RECT  3.800 1.650 3.960 2.060 ;
        RECT  3.550 1.650 3.800 2.050 ;
        RECT  3.030 0.730 3.270 3.490 ;
        RECT  2.410 0.730 3.030 0.970 ;
        RECT  2.250 1.330 2.490 4.180 ;
        RECT  1.120 3.030 2.250 3.270 ;
        RECT  0.720 3.030 1.120 4.010 ;
        RECT  0.500 1.090 0.760 1.490 ;
        RECT  0.500 3.030 0.720 3.270 ;
        RECT  0.260 1.090 0.500 3.270 ;
    END
END DFFSHQX4

MACRO DFFSHQX2
    CLASS CORE ;
    FOREIGN DFFSHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSHQXL ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.190 2.410 4.270 2.870 ;
        RECT  4.270 2.400 4.820 2.870 ;
        RECT  4.820 2.390 5.080 2.870 ;
        RECT  5.080 2.630 5.350 2.870 ;
        RECT  5.350 2.630 5.590 4.350 ;
        RECT  5.590 4.110 7.050 4.350 ;
        RECT  7.050 4.080 7.130 4.350 ;
        RECT  7.130 3.650 7.370 4.350 ;
        RECT  7.370 3.650 8.410 3.890 ;
        RECT  8.410 3.650 8.650 4.370 ;
        RECT  8.650 4.060 8.790 4.370 ;
        RECT  8.790 4.130 11.430 4.370 ;
        RECT  11.430 3.860 11.670 4.370 ;
        RECT  11.670 3.860 12.650 4.100 ;
        RECT  12.650 3.760 12.810 4.100 ;
        RECT  12.810 2.270 13.050 4.100 ;
        RECT  13.050 2.270 13.210 2.670 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.060 2.950 14.120 3.210 ;
        RECT  14.120 2.880 14.520 4.380 ;
        RECT  14.520 2.880 14.730 3.220 ;
        RECT  14.730 2.880 14.780 3.120 ;
        RECT  14.610 1.390 14.780 1.790 ;
        RECT  14.780 1.390 15.010 3.120 ;
        RECT  15.010 1.470 15.020 3.120 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.500 1.830 1.920 2.430 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.670 2.200 1.120 2.800 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.270 5.440 ;
        RECT  1.270 4.480 1.670 5.440 ;
        RECT  1.670 4.640 4.100 5.440 ;
        RECT  4.100 4.190 5.080 5.440 ;
        RECT  5.080 4.640 7.700 5.440 ;
        RECT  7.700 4.170 8.100 5.440 ;
        RECT  8.100 4.640 12.180 5.440 ;
        RECT  12.180 4.480 13.320 5.440 ;
        RECT  13.320 4.080 13.330 5.440 ;
        RECT  13.330 3.820 13.730 5.440 ;
        RECT  13.730 4.640 14.840 5.440 ;
        RECT  14.840 4.340 14.850 5.440 ;
        RECT  14.850 4.140 15.250 5.440 ;
        RECT  15.250 4.340 15.260 5.440 ;
        RECT  15.260 4.640 15.840 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.110 0.400 ;
        RECT  1.110 -0.400 1.120 1.430 ;
        RECT  1.120 -0.400 1.520 1.550 ;
        RECT  1.520 -0.400 1.530 1.430 ;
        RECT  1.530 -0.400 3.620 0.400 ;
        RECT  3.620 -0.400 4.020 0.850 ;
        RECT  4.020 -0.400 6.670 0.400 ;
        RECT  6.670 -0.400 6.910 1.310 ;
        RECT  6.910 -0.400 8.110 0.400 ;
        RECT  8.110 -0.400 8.510 1.310 ;
        RECT  8.510 -0.400 11.710 0.400 ;
        RECT  11.710 -0.400 12.110 0.560 ;
        RECT  12.110 -0.400 13.340 0.400 ;
        RECT  13.340 -0.400 13.740 0.560 ;
        RECT  13.740 -0.400 15.840 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.260 2.070 14.500 2.470 ;
        RECT  14.100 2.070 14.260 2.310 ;
        RECT  13.860 0.860 14.100 2.310 ;
        RECT  11.070 0.860 13.860 1.100 ;
        RECT  12.180 2.120 12.370 3.590 ;
        RECT  12.170 1.790 12.180 3.590 ;
        RECT  12.130 1.390 12.170 3.590 ;
        RECT  11.770 1.390 12.130 2.360 ;
        RECT  11.870 3.350 12.130 3.590 ;
        RECT  11.070 2.760 11.850 3.000 ;
        RECT  11.760 1.790 11.770 2.360 ;
        RECT  11.410 1.960 11.760 2.360 ;
        RECT  10.830 0.860 11.070 3.850 ;
        RECT  10.610 0.860 10.830 1.640 ;
        RECT  9.270 3.610 10.830 3.850 ;
        RECT  10.530 0.830 10.610 1.640 ;
        RECT  10.040 3.090 10.550 3.330 ;
        RECT  10.370 0.830 10.530 1.630 ;
        RECT  9.250 0.830 10.370 1.070 ;
        RECT  9.800 1.310 10.040 3.330 ;
        RECT  9.570 1.310 9.800 1.830 ;
        RECT  8.910 3.090 9.800 3.330 ;
        RECT  7.750 1.590 9.570 1.830 ;
        RECT  6.810 2.110 9.490 2.350 ;
        RECT  9.010 0.830 9.250 1.310 ;
        RECT  8.850 0.910 9.010 1.310 ;
        RECT  8.590 3.090 8.910 3.370 ;
        RECT  7.090 3.130 8.590 3.370 ;
        RECT  7.510 0.910 7.750 1.830 ;
        RECT  7.350 0.910 7.510 1.310 ;
        RECT  6.570 1.590 6.810 3.820 ;
        RECT  6.390 1.590 6.570 1.830 ;
        RECT  5.870 3.580 6.570 3.820 ;
        RECT  6.150 1.360 6.390 1.830 ;
        RECT  6.090 2.110 6.330 2.610 ;
        RECT  6.030 1.360 6.150 1.600 ;
        RECT  5.870 2.110 6.090 2.350 ;
        RECT  5.790 0.670 6.030 1.600 ;
        RECT  5.630 1.870 5.870 2.350 ;
        RECT  5.570 0.670 5.790 0.910 ;
        RECT  5.370 1.870 5.630 2.110 ;
        RECT  4.970 1.350 5.370 2.110 ;
        RECT  4.550 0.790 5.020 1.030 ;
        RECT  3.630 1.870 4.970 2.110 ;
        RECT  3.630 3.390 4.830 3.630 ;
        RECT  4.310 0.790 4.550 1.370 ;
        RECT  3.110 1.130 4.310 1.370 ;
        RECT  3.390 1.870 3.630 3.630 ;
        RECT  2.270 4.060 3.190 4.300 ;
        RECT  2.870 0.670 3.110 3.660 ;
        RECT  2.850 0.670 2.870 1.370 ;
        RECT  2.550 3.420 2.870 3.660 ;
        RECT  2.290 0.670 2.850 0.910 ;
        RECT  2.270 1.960 2.470 3.140 ;
        RECT  2.230 1.960 2.270 4.300 ;
        RECT  2.030 2.900 2.230 4.300 ;
        RECT  0.840 3.080 2.030 3.320 ;
        RECT  0.720 3.080 0.840 3.480 ;
        RECT  0.720 1.250 0.750 1.650 ;
        RECT  0.400 1.240 0.720 1.650 ;
        RECT  0.400 3.080 0.720 3.490 ;
        RECT  0.160 1.240 0.400 3.490 ;
        RECT  0.150 1.240 0.160 1.480 ;
        RECT  0.150 3.250 0.160 3.490 ;
    END
END DFFSHQX2

MACRO DFFSHQX1
    CLASS CORE ;
    FOREIGN DFFSHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSHQXL ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.330 2.290 4.570 2.880 ;
        RECT  4.570 2.380 5.080 2.880 ;
        RECT  5.080 2.640 5.300 2.880 ;
        RECT  5.300 2.640 5.540 4.180 ;
        RECT  5.540 3.940 7.160 4.180 ;
        RECT  7.160 3.940 7.400 4.370 ;
        RECT  7.400 4.080 7.470 4.370 ;
        RECT  7.470 4.130 11.010 4.370 ;
        RECT  11.010 4.060 11.150 4.370 ;
        RECT  11.150 3.940 11.380 4.370 ;
        RECT  11.290 1.960 11.380 2.360 ;
        RECT  11.380 1.960 11.390 4.370 ;
        RECT  11.390 1.960 11.620 4.180 ;
        RECT  11.620 1.960 11.690 2.360 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.910 2.770 12.150 3.470 ;
        RECT  12.150 2.770 12.650 3.010 ;
        RECT  12.650 2.660 12.750 3.010 ;
        RECT  12.740 1.830 12.750 2.090 ;
        RECT  12.710 0.850 12.750 1.500 ;
        RECT  12.750 0.850 12.950 3.010 ;
        RECT  12.950 1.260 12.990 3.010 ;
        RECT  12.990 1.830 13.000 2.090 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.490 1.280 1.520 2.200 ;
        RECT  1.520 1.270 1.730 2.200 ;
        RECT  1.730 1.270 1.780 1.530 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.770 2.140 0.860 2.640 ;
        RECT  0.860 2.140 0.900 2.650 ;
        RECT  0.900 2.130 1.210 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.210 5.440 ;
        RECT  1.210 4.480 1.610 5.440 ;
        RECT  1.610 4.640 4.050 5.440 ;
        RECT  4.050 4.110 5.030 5.440 ;
        RECT  5.030 4.640 6.460 5.440 ;
        RECT  6.460 4.480 6.860 5.440 ;
        RECT  6.860 4.640 11.670 5.440 ;
        RECT  11.670 4.480 12.070 5.440 ;
        RECT  12.070 4.640 12.580 5.440 ;
        RECT  12.580 3.490 12.590 5.440 ;
        RECT  12.590 3.290 12.990 5.440 ;
        RECT  12.990 3.490 13.000 5.440 ;
        RECT  13.000 4.640 13.200 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.090 0.400 ;
        RECT  1.090 -0.400 1.490 0.560 ;
        RECT  1.490 -0.400 3.700 0.400 ;
        RECT  3.700 -0.400 3.710 0.730 ;
        RECT  3.710 -0.400 4.110 0.850 ;
        RECT  4.110 -0.400 4.120 0.730 ;
        RECT  4.120 -0.400 6.750 0.400 ;
        RECT  6.750 -0.400 6.990 1.310 ;
        RECT  6.990 -0.400 9.690 0.400 ;
        RECT  9.690 -0.400 10.090 0.560 ;
        RECT  10.090 -0.400 11.410 0.400 ;
        RECT  11.410 -0.400 11.810 0.980 ;
        RECT  11.810 -0.400 13.200 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.130 1.280 12.370 2.480 ;
        RECT  11.130 1.280 12.130 1.520 ;
        RECT  10.890 0.860 11.130 1.520 ;
        RECT  10.770 0.860 10.890 1.100 ;
        RECT  9.970 3.570 10.870 3.810 ;
        RECT  10.370 0.690 10.770 1.100 ;
        RECT  10.150 1.380 10.390 2.710 ;
        RECT  9.870 0.860 10.370 1.100 ;
        RECT  9.970 2.470 10.150 2.710 ;
        RECT  9.730 2.470 9.970 3.810 ;
        RECT  9.630 0.860 9.870 2.190 ;
        RECT  9.410 0.860 9.630 1.100 ;
        RECT  9.450 1.950 9.630 2.190 ;
        RECT  9.210 1.950 9.450 3.130 ;
        RECT  9.120 0.780 9.410 1.100 ;
        RECT  8.220 2.890 9.210 3.130 ;
        RECT  6.730 3.410 9.190 3.650 ;
        RECT  8.350 0.780 9.120 1.020 ;
        RECT  8.270 1.380 9.050 1.620 ;
        RECT  8.030 1.380 8.270 2.370 ;
        RECT  7.810 2.130 8.030 2.370 ;
        RECT  7.570 2.130 7.810 2.610 ;
        RECT  7.510 0.910 7.750 1.840 ;
        RECT  7.250 2.890 7.740 3.130 ;
        RECT  7.250 1.600 7.510 1.840 ;
        RECT  7.010 1.600 7.250 3.130 ;
        RECT  6.490 1.590 6.730 3.650 ;
        RECT  6.470 1.590 6.490 1.830 ;
        RECT  6.370 3.390 6.490 3.650 ;
        RECT  6.230 1.360 6.470 1.830 ;
        RECT  5.870 3.390 6.370 3.630 ;
        RECT  6.010 2.110 6.250 2.670 ;
        RECT  6.110 1.360 6.230 1.600 ;
        RECT  5.870 0.670 6.110 1.600 ;
        RECT  5.690 2.110 6.010 2.350 ;
        RECT  5.650 0.670 5.870 0.910 ;
        RECT  5.450 1.840 5.690 2.350 ;
        RECT  5.210 1.340 5.450 2.080 ;
        RECT  4.630 0.770 5.250 1.010 ;
        RECT  5.050 1.340 5.210 2.000 ;
        RECT  4.050 1.760 5.050 2.000 ;
        RECT  4.050 3.390 4.830 3.630 ;
        RECT  4.390 0.770 4.630 1.370 ;
        RECT  3.290 1.130 4.390 1.370 ;
        RECT  3.810 1.760 4.050 3.630 ;
        RECT  3.570 1.760 3.810 2.160 ;
        RECT  3.290 2.440 3.530 4.050 ;
        RECT  3.280 0.670 3.290 1.370 ;
        RECT  3.280 2.440 3.290 2.680 ;
        RECT  2.550 3.810 3.290 4.050 ;
        RECT  3.040 0.670 3.280 2.680 ;
        RECT  2.290 0.670 3.040 0.910 ;
        RECT  2.770 3.130 3.010 3.530 ;
        RECT  2.450 3.290 2.770 3.530 ;
        RECT  2.210 1.810 2.450 3.530 ;
        RECT  0.780 3.290 2.210 3.530 ;
        RECT  0.480 3.290 0.780 3.780 ;
        RECT  0.480 1.230 0.670 1.630 ;
        RECT  0.240 1.230 0.480 3.780 ;
    END
END DFFSHQX1

MACRO DFFSXL
    CLASS CORE ;
    FOREIGN DFFSXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.440 4.070 9.450 4.330 ;
        RECT  9.450 4.060 9.700 4.330 ;
        RECT  9.700 4.060 9.840 4.300 ;
        RECT  9.840 3.740 10.080 4.300 ;
        RECT  10.080 3.740 10.240 4.140 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.170 3.520 11.420 3.950 ;
        RECT  11.420 3.510 11.570 3.950 ;
        RECT  11.230 0.690 11.630 1.100 ;
        RECT  11.570 3.510 11.680 3.770 ;
        RECT  11.630 0.860 11.990 1.100 ;
        RECT  11.680 3.520 12.130 3.760 ;
        RECT  11.990 0.860 12.130 1.280 ;
        RECT  12.130 0.860 12.370 3.760 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.650 3.160 12.700 3.560 ;
        RECT  12.700 1.280 13.000 3.570 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.330 1.280 1.520 2.240 ;
        RECT  1.520 1.270 1.570 2.240 ;
        RECT  1.570 1.270 1.780 1.530 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.560 0.800 3.200 ;
        RECT  0.800 2.550 0.860 3.200 ;
        RECT  0.860 2.550 1.120 3.210 ;
        RECT  1.120 2.550 1.130 2.970 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.090 5.440 ;
        RECT  1.090 4.480 1.490 5.440 ;
        RECT  1.490 4.640 3.490 5.440 ;
        RECT  3.490 4.480 3.890 5.440 ;
        RECT  3.890 4.640 5.020 5.440 ;
        RECT  5.020 4.310 5.030 5.440 ;
        RECT  5.030 4.190 5.430 5.440 ;
        RECT  5.430 4.310 5.440 5.440 ;
        RECT  5.440 4.640 6.340 5.440 ;
        RECT  6.340 4.310 6.350 5.440 ;
        RECT  6.350 4.190 6.750 5.440 ;
        RECT  6.750 4.310 6.760 5.440 ;
        RECT  6.760 4.640 8.640 5.440 ;
        RECT  8.640 4.210 8.650 5.440 ;
        RECT  8.650 4.010 9.050 5.440 ;
        RECT  9.050 4.210 9.060 5.440 ;
        RECT  9.060 4.640 10.490 5.440 ;
        RECT  10.490 3.730 10.730 5.440 ;
        RECT  10.730 4.640 11.960 5.440 ;
        RECT  11.960 4.480 12.360 5.440 ;
        RECT  12.360 4.640 13.200 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.910 0.400 ;
        RECT  0.910 -0.400 1.310 0.560 ;
        RECT  1.310 -0.400 3.600 0.400 ;
        RECT  3.600 -0.400 3.610 0.750 ;
        RECT  3.610 -0.400 4.010 0.870 ;
        RECT  4.010 -0.400 4.020 0.750 ;
        RECT  4.020 -0.400 6.000 0.400 ;
        RECT  6.000 -0.400 6.010 0.730 ;
        RECT  6.010 -0.400 6.410 0.850 ;
        RECT  6.410 -0.400 6.420 0.730 ;
        RECT  6.420 -0.400 8.270 0.400 ;
        RECT  8.270 -0.400 8.670 0.560 ;
        RECT  8.670 -0.400 10.340 0.400 ;
        RECT  10.340 -0.400 10.350 0.850 ;
        RECT  10.350 -0.400 10.750 1.050 ;
        RECT  10.750 -0.400 10.760 0.850 ;
        RECT  10.760 -0.400 11.970 0.400 ;
        RECT  11.970 -0.400 12.370 0.560 ;
        RECT  12.370 -0.400 13.200 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  11.640 1.960 11.850 2.370 ;
        RECT  11.630 1.500 11.640 2.370 ;
        RECT  11.390 1.380 11.630 3.210 ;
        RECT  11.380 1.380 11.390 2.110 ;
        RECT  11.230 2.810 11.390 3.210 ;
        RECT  11.230 1.380 11.380 1.780 ;
        RECT  10.790 2.020 10.950 2.420 ;
        RECT  10.550 1.570 10.790 3.210 ;
        RECT  9.410 1.570 10.550 1.810 ;
        RECT  9.930 2.970 10.550 3.210 ;
        RECT  9.530 2.970 9.930 3.370 ;
        RECT  9.230 2.290 9.630 2.690 ;
        RECT  9.010 1.220 9.410 1.810 ;
        RECT  8.230 2.370 9.230 2.610 ;
        RECT  8.750 1.570 9.010 1.810 ;
        RECT  8.510 1.570 8.750 1.970 ;
        RECT  7.990 1.490 8.230 4.370 ;
        RECT  7.470 1.490 7.990 1.730 ;
        RECT  7.470 2.730 7.710 3.910 ;
        RECT  7.230 1.330 7.470 1.730 ;
        RECT  5.950 3.670 7.470 3.910 ;
        RECT  6.950 2.010 7.250 2.410 ;
        RECT  6.710 1.240 6.950 3.390 ;
        RECT  5.570 1.240 6.710 1.480 ;
        RECT  5.910 3.150 6.710 3.390 ;
        RECT  6.190 2.020 6.430 2.420 ;
        RECT  5.520 2.100 6.190 2.340 ;
        RECT  5.710 3.670 5.950 4.070 ;
        RECT  3.210 3.670 5.710 3.910 ;
        RECT  5.330 0.670 5.570 1.480 ;
        RECT  5.280 1.760 5.520 3.400 ;
        RECT  4.560 0.670 5.330 0.910 ;
        RECT  5.050 1.760 5.280 2.000 ;
        RECT  3.570 3.160 5.280 3.400 ;
        RECT  4.810 1.430 5.050 2.000 ;
        RECT  4.750 2.370 4.990 2.770 ;
        RECT  4.280 2.370 4.750 2.610 ;
        RECT  4.040 1.210 4.280 2.610 ;
        RECT  2.890 1.210 4.040 1.450 ;
        RECT  3.330 2.160 3.570 3.400 ;
        RECT  2.970 3.670 3.210 4.140 ;
        RECT  2.170 3.900 2.970 4.140 ;
        RECT  2.690 1.210 2.890 2.910 ;
        RECT  2.670 1.210 2.690 3.500 ;
        RECT  2.650 1.050 2.670 3.500 ;
        RECT  2.270 1.050 2.650 1.450 ;
        RECT  2.450 2.670 2.650 3.500 ;
        RECT  2.170 1.810 2.370 2.050 ;
        RECT  1.930 1.810 2.170 4.140 ;
        RECT  0.570 3.900 1.930 4.140 ;
        RECT  0.400 1.270 0.570 1.670 ;
        RECT  0.400 3.490 0.570 4.140 ;
        RECT  0.330 1.270 0.400 4.140 ;
        RECT  0.160 1.270 0.330 3.890 ;
    END
END DFFSXL

MACRO DFFSX4
    CLASS CORE ;
    FOREIGN DFFSX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSXL ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.070 4.060 4.690 4.380 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.680 1.580 15.690 2.730 ;
        RECT  15.690 1.380 15.700 2.730 ;
        RECT  15.700 1.380 15.710 2.950 ;
        RECT  15.710 1.380 15.950 3.150 ;
        RECT  15.950 1.380 16.090 3.220 ;
        RECT  16.090 1.580 16.100 3.220 ;
        RECT  16.100 1.820 16.390 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.220 1.380 17.250 2.730 ;
        RECT  17.250 1.380 17.270 3.150 ;
        RECT  17.270 1.380 17.710 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.240 1.560 1.430 1.960 ;
        RECT  1.430 1.270 1.780 1.970 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.770 2.290 1.460 2.690 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.130 5.440 ;
        RECT  1.130 4.480 1.530 5.440 ;
        RECT  1.530 4.640 3.560 5.440 ;
        RECT  3.560 4.170 3.800 5.440 ;
        RECT  3.800 4.640 5.010 5.440 ;
        RECT  5.010 4.310 5.020 5.440 ;
        RECT  5.020 4.110 5.420 5.440 ;
        RECT  5.420 4.310 5.430 5.440 ;
        RECT  5.430 4.640 6.350 5.440 ;
        RECT  6.350 4.310 6.360 5.440 ;
        RECT  6.360 4.110 6.760 5.440 ;
        RECT  6.760 4.310 6.770 5.440 ;
        RECT  6.770 4.640 8.900 5.440 ;
        RECT  8.900 3.630 9.300 5.440 ;
        RECT  9.300 4.640 10.730 5.440 ;
        RECT  10.730 4.010 11.130 5.440 ;
        RECT  11.130 4.640 12.120 5.440 ;
        RECT  12.120 3.660 12.130 5.440 ;
        RECT  12.130 3.460 12.530 5.440 ;
        RECT  12.530 3.660 12.540 5.440 ;
        RECT  12.540 4.640 13.350 5.440 ;
        RECT  13.350 4.630 13.530 5.440 ;
        RECT  13.530 3.500 13.930 5.440 ;
        RECT  13.930 4.640 15.100 5.440 ;
        RECT  15.100 4.010 15.500 5.440 ;
        RECT  15.500 4.640 16.480 5.440 ;
        RECT  16.480 4.210 16.490 5.440 ;
        RECT  16.490 4.010 16.890 5.440 ;
        RECT  16.890 4.210 16.900 5.440 ;
        RECT  16.900 4.640 17.920 5.440 ;
        RECT  17.920 4.010 18.320 5.440 ;
        RECT  18.320 4.640 18.480 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.140 0.400 ;
        RECT  1.140 -0.400 1.540 0.560 ;
        RECT  1.540 -0.400 3.590 0.400 ;
        RECT  3.590 -0.400 3.600 1.000 ;
        RECT  3.600 -0.400 4.000 1.120 ;
        RECT  4.000 -0.400 4.010 1.000 ;
        RECT  4.010 -0.400 6.490 0.400 ;
        RECT  6.490 -0.400 6.500 1.010 ;
        RECT  6.500 -0.400 6.900 1.130 ;
        RECT  6.900 -0.400 6.910 1.010 ;
        RECT  6.910 -0.400 9.130 0.400 ;
        RECT  9.130 -0.400 9.140 0.840 ;
        RECT  9.140 -0.400 9.540 0.960 ;
        RECT  9.540 -0.400 9.550 0.840 ;
        RECT  9.550 -0.400 10.970 0.400 ;
        RECT  10.970 -0.400 11.370 0.560 ;
        RECT  11.370 -0.400 13.520 0.400 ;
        RECT  13.520 -0.400 13.530 1.020 ;
        RECT  13.530 -0.400 13.930 1.220 ;
        RECT  13.930 -0.400 13.940 1.020 ;
        RECT  13.940 -0.400 15.070 0.400 ;
        RECT  15.070 -0.400 15.080 0.900 ;
        RECT  15.080 -0.400 15.480 1.100 ;
        RECT  15.480 -0.400 15.490 0.900 ;
        RECT  15.490 -0.400 16.460 0.400 ;
        RECT  16.460 -0.400 16.470 0.900 ;
        RECT  16.470 -0.400 16.870 1.100 ;
        RECT  16.870 -0.400 16.880 0.900 ;
        RECT  16.880 -0.400 17.890 0.400 ;
        RECT  17.890 -0.400 17.900 0.900 ;
        RECT  17.900 -0.400 18.300 1.100 ;
        RECT  18.300 -0.400 18.310 0.900 ;
        RECT  18.310 -0.400 18.480 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  17.990 2.150 18.230 3.730 ;
        RECT  15.230 3.490 17.990 3.730 ;
        RECT  14.990 1.390 15.230 3.730 ;
        RECT  14.680 1.390 14.990 1.630 ;
        RECT  14.250 2.750 14.990 3.150 ;
        RECT  14.470 2.050 14.710 2.450 ;
        RECT  14.280 1.200 14.680 1.630 ;
        RECT  13.400 2.050 14.470 2.440 ;
        RECT  13.160 1.500 13.400 2.440 ;
        RECT  13.140 2.780 13.200 3.180 ;
        RECT  12.650 1.500 13.160 1.740 ;
        RECT  13.140 2.200 13.160 2.440 ;
        RECT  12.900 2.200 13.140 3.180 ;
        RECT  12.800 2.780 12.900 3.180 ;
        RECT  11.670 2.860 12.800 3.100 ;
        RECT  12.250 1.210 12.650 1.740 ;
        RECT  12.110 2.180 12.510 2.580 ;
        RECT  11.080 1.500 12.250 1.740 ;
        RECT  10.200 2.340 12.110 2.580 ;
        RECT  11.430 2.860 11.670 3.730 ;
        RECT  11.400 2.860 11.430 3.100 ;
        RECT  10.490 3.490 11.430 3.730 ;
        RECT  10.840 1.500 11.080 2.060 ;
        RECT  10.680 1.820 10.840 2.060 ;
        RECT  10.250 3.490 10.490 4.070 ;
        RECT  9.960 1.240 10.200 3.200 ;
        RECT  9.660 1.240 9.960 1.700 ;
        RECT  7.960 2.960 9.960 3.200 ;
        RECT  9.440 2.170 9.680 2.570 ;
        RECT  8.260 1.240 9.660 1.480 ;
        RECT  8.520 2.250 9.440 2.490 ;
        RECT  8.280 1.760 8.520 2.490 ;
        RECT  6.940 1.760 8.280 2.000 ;
        RECT  8.020 1.130 8.260 1.480 ;
        RECT  7.860 1.130 8.020 1.370 ;
        RECT  7.720 2.960 7.960 3.470 ;
        RECT  7.440 2.360 7.800 2.600 ;
        RECT  7.200 2.360 7.440 3.830 ;
        RECT  5.940 3.590 7.200 3.830 ;
        RECT  6.920 1.410 6.940 2.000 ;
        RECT  6.680 1.410 6.920 3.270 ;
        RECT  5.940 1.410 6.680 1.650 ;
        RECT  5.840 3.030 6.680 3.270 ;
        RECT  6.160 2.240 6.400 2.640 ;
        RECT  5.560 2.320 6.160 2.560 ;
        RECT  5.700 0.670 5.940 1.650 ;
        RECT  5.700 3.550 5.940 4.130 ;
        RECT  5.560 0.670 5.700 1.070 ;
        RECT  3.280 3.550 5.700 3.790 ;
        RECT  5.320 1.930 5.560 3.270 ;
        RECT  5.200 1.930 5.320 2.170 ;
        RECT  4.100 3.030 5.320 3.270 ;
        RECT  4.960 0.930 5.200 2.170 ;
        RECT  4.630 2.450 5.040 2.690 ;
        RECT  4.390 1.400 4.630 2.690 ;
        RECT  2.900 1.400 4.390 1.640 ;
        RECT  3.860 2.090 4.100 3.270 ;
        RECT  3.780 2.090 3.860 2.330 ;
        RECT  3.540 1.930 3.780 2.330 ;
        RECT  3.040 3.550 3.280 4.290 ;
        RECT  2.240 4.050 3.040 4.290 ;
        RECT  2.760 1.400 2.900 3.130 ;
        RECT  2.660 1.400 2.760 3.760 ;
        RECT  2.420 1.000 2.660 1.640 ;
        RECT  2.520 2.890 2.660 3.760 ;
        RECT  2.260 1.000 2.420 1.400 ;
        RECT  2.240 1.990 2.380 2.610 ;
        RECT  2.140 1.990 2.240 4.290 ;
        RECT  2.000 2.370 2.140 4.290 ;
        RECT  0.670 3.870 2.000 4.110 ;
        RECT  0.500 0.940 0.670 1.340 ;
        RECT  0.500 2.970 0.670 4.110 ;
        RECT  0.430 0.940 0.500 4.110 ;
        RECT  0.260 0.940 0.430 3.370 ;
    END
END DFFSX4

MACRO DFFSX2
    CLASS CORE ;
    FOREIGN DFFSX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.520 2.090 ;
        RECT  3.520 1.830 3.760 2.100 ;
        RECT  3.760 1.860 3.920 2.100 ;
        RECT  3.920 1.860 4.160 2.400 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.850 2.750 11.990 3.150 ;
        RECT  11.990 2.380 12.080 3.150 ;
        RECT  11.730 0.710 12.080 0.950 ;
        RECT  12.080 0.710 12.320 3.150 ;
        RECT  12.320 2.390 12.330 3.150 ;
        RECT  12.330 2.390 12.340 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.740 1.260 13.290 1.540 ;
        RECT  13.290 2.760 13.370 3.900 ;
        RECT  13.290 1.260 13.370 1.670 ;
        RECT  13.370 1.260 13.690 3.900 ;
        RECT  13.690 1.260 13.700 2.980 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.200 1.870 1.280 2.110 ;
        RECT  1.280 1.280 1.520 2.110 ;
        RECT  1.520 1.870 1.600 2.110 ;
        RECT  1.520 1.270 1.780 1.530 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.380 1.210 2.910 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.920 5.440 ;
        RECT  0.920 4.480 1.320 5.440 ;
        RECT  1.320 4.640 3.350 5.440 ;
        RECT  3.350 4.480 3.750 5.440 ;
        RECT  3.750 4.640 4.870 5.440 ;
        RECT  4.870 4.310 4.880 5.440 ;
        RECT  4.880 4.190 5.280 5.440 ;
        RECT  5.280 4.310 5.290 5.440 ;
        RECT  5.290 4.640 6.270 5.440 ;
        RECT  6.270 4.220 6.280 5.440 ;
        RECT  6.280 4.020 6.680 5.440 ;
        RECT  6.680 4.220 6.690 5.440 ;
        RECT  6.690 4.640 8.770 5.440 ;
        RECT  8.770 4.010 9.010 5.440 ;
        RECT  9.010 4.640 10.270 5.440 ;
        RECT  10.270 3.520 10.670 5.440 ;
        RECT  10.670 4.640 12.530 5.440 ;
        RECT  12.530 4.090 12.930 5.440 ;
        RECT  12.930 4.640 13.860 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.830 0.400 ;
        RECT  0.830 -0.400 1.230 0.560 ;
        RECT  1.230 -0.400 3.550 0.400 ;
        RECT  3.550 -0.400 3.560 0.910 ;
        RECT  3.560 -0.400 3.960 1.030 ;
        RECT  3.960 -0.400 3.970 0.910 ;
        RECT  3.970 -0.400 6.020 0.400 ;
        RECT  6.020 -0.400 6.260 1.110 ;
        RECT  6.260 -0.400 8.560 0.400 ;
        RECT  8.560 -0.400 8.960 0.960 ;
        RECT  8.960 -0.400 10.530 0.400 ;
        RECT  10.530 -0.400 10.930 0.560 ;
        RECT  10.930 -0.400 12.610 0.400 ;
        RECT  12.610 -0.400 12.850 0.930 ;
        RECT  12.850 -0.400 13.860 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.940 1.990 13.090 2.390 ;
        RECT  12.700 1.990 12.940 3.740 ;
        RECT  11.570 3.500 12.700 3.740 ;
        RECT  11.570 1.470 11.590 1.710 ;
        RECT  11.430 1.470 11.570 3.740 ;
        RECT  11.330 1.470 11.430 3.900 ;
        RECT  11.190 1.470 11.330 1.710 ;
        RECT  11.030 3.500 11.330 3.900 ;
        RECT  10.910 2.020 11.050 2.450 ;
        RECT  10.670 1.500 10.910 3.220 ;
        RECT  9.650 1.500 10.670 1.740 ;
        RECT  9.910 2.980 10.670 3.220 ;
        RECT  9.750 2.980 9.910 3.380 ;
        RECT  9.510 2.980 9.750 3.730 ;
        RECT  9.250 1.240 9.650 1.740 ;
        RECT  8.470 3.490 9.510 3.730 ;
        RECT  9.090 2.100 9.490 2.500 ;
        RECT  8.260 1.240 9.250 1.480 ;
        RECT  7.880 2.180 9.090 2.420 ;
        RECT  8.230 3.490 8.470 4.070 ;
        RECT  8.070 3.670 8.230 4.070 ;
        RECT  7.640 1.300 7.880 3.330 ;
        RECT  7.360 3.950 7.720 4.190 ;
        RECT  7.540 1.300 7.640 1.540 ;
        RECT  7.300 1.140 7.540 1.540 ;
        RECT  7.020 1.820 7.360 2.060 ;
        RECT  7.120 3.500 7.360 4.190 ;
        RECT  6.000 3.500 7.120 3.740 ;
        RECT  6.780 1.410 7.020 3.120 ;
        RECT  5.740 1.410 6.780 1.650 ;
        RECT  5.760 2.880 6.780 3.120 ;
        RECT  6.260 2.150 6.500 2.550 ;
        RECT  5.480 2.230 6.260 2.470 ;
        RECT  5.800 3.500 6.000 3.920 ;
        RECT  5.760 3.500 5.800 4.080 ;
        RECT  5.560 3.670 5.760 4.080 ;
        RECT  5.500 0.670 5.740 1.650 ;
        RECT  3.060 3.670 5.560 3.910 ;
        RECT  4.490 0.670 5.500 0.910 ;
        RECT  5.240 1.930 5.480 3.390 ;
        RECT  5.220 1.930 5.240 2.170 ;
        RECT  3.400 3.150 5.240 3.390 ;
        RECT  4.980 1.440 5.220 2.170 ;
        RECT  4.700 2.510 4.920 2.750 ;
        RECT  4.460 1.310 4.700 2.750 ;
        RECT  2.880 1.310 4.460 1.550 ;
        RECT  3.160 2.410 3.400 3.390 ;
        RECT  2.820 3.670 3.060 4.210 ;
        RECT  2.640 0.850 2.880 3.300 ;
        RECT  2.020 3.970 2.820 4.210 ;
        RECT  2.220 0.850 2.640 1.250 ;
        RECT  2.540 3.060 2.640 3.300 ;
        RECT  2.300 3.060 2.540 3.580 ;
        RECT  2.020 1.810 2.240 2.780 ;
        RECT  2.000 1.810 2.020 4.210 ;
        RECT  1.780 2.540 2.000 4.210 ;
        RECT  0.570 3.350 1.780 3.590 ;
        RECT  0.400 1.220 0.570 1.620 ;
        RECT  0.400 3.190 0.570 3.590 ;
        RECT  0.160 1.220 0.400 3.590 ;
    END
END DFFSX2

MACRO DFFSX1
    CLASS CORE ;
    FOREIGN DFFSX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFSXL ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.440 4.070 9.450 4.330 ;
        RECT  9.450 3.900 9.700 4.330 ;
        RECT  9.700 3.900 9.780 4.140 ;
        RECT  9.780 3.740 10.020 4.140 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  10.990 0.670 11.250 0.910 ;
        RECT  11.040 3.650 11.420 4.050 ;
        RECT  11.250 0.670 11.490 1.100 ;
        RECT  11.420 3.500 11.670 4.050 ;
        RECT  11.670 3.500 11.680 3.770 ;
        RECT  11.680 3.500 11.880 3.760 ;
        RECT  11.490 0.860 11.880 1.100 ;
        RECT  11.880 0.860 12.120 3.760 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.520 2.840 12.650 3.240 ;
        RECT  12.470 1.220 12.650 1.620 ;
        RECT  12.650 1.220 12.740 1.820 ;
        RECT  12.650 2.660 12.750 3.240 ;
        RECT  12.740 1.220 12.750 2.090 ;
        RECT  12.750 1.220 12.760 3.240 ;
        RECT  12.760 1.220 12.980 3.080 ;
        RECT  12.980 1.830 12.990 3.080 ;
        RECT  12.990 1.830 13.000 2.090 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.220 1.670 1.780 2.090 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.690 0.790 3.200 ;
        RECT  0.790 2.680 0.860 3.200 ;
        RECT  0.860 2.680 1.120 3.210 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.010 5.440 ;
        RECT  1.010 4.480 1.410 5.440 ;
        RECT  1.410 4.640 3.560 5.440 ;
        RECT  3.560 4.480 3.960 5.440 ;
        RECT  3.960 4.640 4.980 5.440 ;
        RECT  4.980 4.210 4.990 5.440 ;
        RECT  4.990 4.090 5.390 5.440 ;
        RECT  5.390 4.210 5.400 5.440 ;
        RECT  5.400 4.640 6.320 5.440 ;
        RECT  6.320 4.110 6.560 5.440 ;
        RECT  6.560 4.640 8.630 5.440 ;
        RECT  8.630 4.310 8.640 5.440 ;
        RECT  8.640 4.110 9.040 5.440 ;
        RECT  9.040 4.310 9.050 5.440 ;
        RECT  9.050 4.640 10.300 5.440 ;
        RECT  10.300 3.080 10.540 5.440 ;
        RECT  10.540 4.640 11.830 5.440 ;
        RECT  11.830 4.480 12.230 5.440 ;
        RECT  12.230 4.640 13.200 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.870 0.400 ;
        RECT  0.870 -0.400 1.270 0.560 ;
        RECT  1.270 -0.400 3.580 0.400 ;
        RECT  3.580 -0.400 3.590 0.880 ;
        RECT  3.590 -0.400 3.990 1.000 ;
        RECT  3.990 -0.400 4.000 0.880 ;
        RECT  4.000 -0.400 5.830 0.400 ;
        RECT  5.830 -0.400 6.070 0.950 ;
        RECT  6.070 -0.400 8.210 0.400 ;
        RECT  8.210 -0.400 8.610 0.560 ;
        RECT  8.610 -0.400 10.220 0.400 ;
        RECT  10.220 -0.400 10.230 0.670 ;
        RECT  10.230 -0.400 10.630 0.870 ;
        RECT  10.630 -0.400 10.640 0.670 ;
        RECT  10.640 -0.400 11.770 0.400 ;
        RECT  11.770 -0.400 12.170 0.560 ;
        RECT  12.170 -0.400 13.200 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  11.500 2.080 11.580 2.480 ;
        RECT  11.260 1.380 11.500 3.230 ;
        RECT  11.050 1.380 11.260 1.780 ;
        RECT  11.100 2.990 11.260 3.230 ;
        RECT  10.420 2.110 10.820 2.510 ;
        RECT  9.860 2.190 10.420 2.430 ;
        RECT  9.620 1.630 9.860 3.430 ;
        RECT  9.350 1.630 9.620 1.870 ;
        RECT  9.460 3.030 9.620 3.430 ;
        RECT  8.950 1.160 9.350 1.870 ;
        RECT  9.080 2.350 9.320 2.750 ;
        RECT  7.980 2.430 9.080 2.670 ;
        RECT  8.700 1.630 8.950 1.870 ;
        RECT  8.300 1.630 8.700 2.030 ;
        RECT  7.840 1.230 7.980 3.760 ;
        RECT  7.740 1.230 7.840 3.920 ;
        RECT  7.090 1.230 7.740 1.470 ;
        RECT  7.600 3.520 7.740 3.920 ;
        RECT  7.320 2.520 7.460 2.920 ;
        RECT  7.080 2.520 7.320 3.810 ;
        RECT  6.800 1.840 7.180 2.080 ;
        RECT  3.420 3.570 7.080 3.810 ;
        RECT  6.560 1.230 6.800 2.920 ;
        RECT  5.550 1.230 6.560 1.470 ;
        RECT  6.290 2.680 6.560 2.920 ;
        RECT  6.050 2.680 6.290 3.180 ;
        RECT  6.040 1.750 6.280 2.150 ;
        RECT  5.750 1.830 6.040 2.070 ;
        RECT  5.510 1.830 5.750 3.290 ;
        RECT  5.310 0.670 5.550 1.470 ;
        RECT  5.030 1.830 5.510 2.070 ;
        RECT  3.650 3.050 5.510 3.290 ;
        RECT  4.300 0.670 5.310 0.910 ;
        RECT  4.790 1.370 5.030 2.070 ;
        RECT  4.650 2.350 4.890 2.770 ;
        RECT  4.330 2.350 4.650 2.590 ;
        RECT  4.090 1.280 4.330 2.590 ;
        RECT  2.900 1.280 4.090 1.520 ;
        RECT  3.410 2.370 3.650 3.290 ;
        RECT  3.180 3.570 3.420 4.160 ;
        RECT  3.250 2.370 3.410 2.770 ;
        RECT  2.230 3.920 3.180 4.160 ;
        RECT  2.660 0.850 2.900 3.640 ;
        RECT  2.250 0.850 2.660 1.250 ;
        RECT  2.510 3.240 2.660 3.640 ;
        RECT  2.230 1.530 2.380 2.610 ;
        RECT  2.140 1.530 2.230 4.160 ;
        RECT  1.990 2.370 2.140 4.160 ;
        RECT  0.570 3.570 1.990 3.810 ;
        RECT  0.400 1.140 0.570 1.540 ;
        RECT  0.400 3.490 0.570 3.890 ;
        RECT  0.160 1.140 0.400 3.890 ;
    END
END DFFSX1

MACRO DFFRHQXL
    CLASS CORE ;
    FOREIGN DFFRHQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  11.850 2.910 12.430 3.260 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.710 1.000 12.950 1.400 ;
        RECT  13.280 3.690 13.350 4.090 ;
        RECT  13.350 3.040 13.400 4.100 ;
        RECT  13.400 2.950 13.450 4.100 ;
        RECT  12.950 1.160 13.450 1.400 ;
        RECT  13.450 1.160 13.690 4.100 ;
        RECT  13.690 3.040 13.700 4.100 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.630 2.090 ;
        RECT  1.630 1.830 1.780 2.460 ;
        RECT  1.780 1.840 1.870 2.460 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.770 2.210 1.170 2.730 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.300 5.440 ;
        RECT  1.300 3.650 1.310 5.440 ;
        RECT  1.310 3.530 1.710 5.440 ;
        RECT  1.710 3.650 1.720 5.440 ;
        RECT  1.720 4.640 3.920 5.440 ;
        RECT  3.920 4.280 3.930 5.440 ;
        RECT  3.930 4.160 4.330 5.440 ;
        RECT  4.330 4.280 4.340 5.440 ;
        RECT  4.340 4.640 7.330 5.440 ;
        RECT  7.330 4.480 7.730 5.440 ;
        RECT  7.730 4.640 9.920 5.440 ;
        RECT  9.920 4.480 10.320 5.440 ;
        RECT  11.130 3.180 11.530 3.770 ;
        RECT  10.320 4.640 12.060 5.440 ;
        RECT  11.530 3.530 12.060 3.770 ;
        RECT  12.060 3.530 12.300 5.440 ;
        RECT  12.300 3.740 12.460 5.440 ;
        RECT  12.460 4.640 13.860 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.360 0.400 ;
        RECT  1.360 -0.400 1.370 1.430 ;
        RECT  1.370 -0.400 1.770 1.550 ;
        RECT  1.770 -0.400 1.780 1.430 ;
        RECT  1.780 -0.400 3.900 0.400 ;
        RECT  3.900 -0.400 4.060 1.170 ;
        RECT  4.060 -0.400 4.300 1.440 ;
        RECT  4.300 1.200 5.440 1.440 ;
        RECT  5.440 1.190 5.450 1.540 ;
        RECT  5.450 1.190 5.850 1.830 ;
        RECT  5.850 1.190 5.860 1.540 ;
        RECT  4.300 -0.400 6.650 0.400 ;
        RECT  6.650 -0.400 7.070 1.170 ;
        RECT  7.070 -0.400 9.570 0.400 ;
        RECT  9.570 -0.400 9.970 0.560 ;
        RECT  9.970 -0.400 11.180 0.400 ;
        RECT  11.180 -0.400 12.160 0.560 ;
        RECT  12.160 -0.400 13.300 0.400 ;
        RECT  13.300 -0.400 13.700 0.560 ;
        RECT  13.700 -0.400 13.860 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.930 1.680 13.170 2.080 ;
        RECT  12.700 2.400 12.940 2.810 ;
        RECT  12.430 1.760 12.930 2.000 ;
        RECT  11.730 2.400 12.700 2.640 ;
        RECT  12.190 0.860 12.430 2.000 ;
        RECT  10.320 0.860 12.190 1.100 ;
        RECT  11.490 1.660 11.730 2.640 ;
        RECT  10.850 4.090 11.580 4.330 ;
        RECT  11.330 1.660 11.490 1.900 ;
        RECT  10.850 2.400 11.490 2.640 ;
        RECT  10.610 2.400 10.850 4.330 ;
        RECT  10.150 1.470 10.670 1.710 ;
        RECT  5.810 3.940 10.610 4.180 ;
        RECT  9.920 0.860 10.320 1.150 ;
        RECT  10.150 3.210 10.310 3.610 ;
        RECT  9.910 1.470 10.150 3.610 ;
        RECT  9.570 0.860 9.920 1.100 ;
        RECT  9.610 2.680 9.910 2.920 ;
        RECT  9.330 0.860 9.570 2.360 ;
        RECT  8.550 0.860 9.330 1.110 ;
        RECT  9.210 2.120 9.330 2.360 ;
        RECT  8.970 2.120 9.210 3.660 ;
        RECT  8.590 3.420 8.970 3.660 ;
        RECT  8.690 1.600 8.950 1.840 ;
        RECT  8.450 1.600 8.690 3.140 ;
        RECT  8.310 0.860 8.550 1.320 ;
        RECT  8.170 3.420 8.230 3.660 ;
        RECT  8.030 1.590 8.170 3.660 ;
        RECT  7.930 1.060 8.030 3.660 ;
        RECT  7.790 1.060 7.930 1.830 ;
        RECT  7.830 3.420 7.930 3.660 ;
        RECT  7.460 1.060 7.790 1.300 ;
        RECT  7.510 2.300 7.650 2.700 ;
        RECT  7.270 1.580 7.510 3.660 ;
        RECT  6.380 1.580 7.270 1.820 ;
        RECT  6.430 3.420 7.270 3.660 ;
        RECT  6.690 2.170 6.930 2.600 ;
        RECT  5.130 2.170 6.690 2.410 ;
        RECT  6.140 0.680 6.380 1.820 ;
        RECT  4.590 0.680 6.140 0.920 ;
        RECT  5.570 2.690 5.810 4.180 ;
        RECT  5.410 2.690 5.570 2.930 ;
        RECT  4.970 2.030 5.130 3.550 ;
        RECT  4.890 1.720 4.970 3.550 ;
        RECT  4.570 1.720 4.890 2.270 ;
        RECT  4.770 3.310 4.890 3.550 ;
        RECT  4.530 3.310 4.770 3.710 ;
        RECT  4.350 2.550 4.590 2.950 ;
        RECT  3.870 2.030 4.570 2.270 ;
        RECT  3.290 2.710 4.350 2.950 ;
        RECT  3.630 2.000 3.870 2.400 ;
        RECT  3.050 0.670 3.290 3.320 ;
        RECT  2.390 4.100 3.290 4.340 ;
        RECT  2.570 0.670 3.050 0.910 ;
        RECT  2.910 3.080 3.050 3.320 ;
        RECT  2.670 3.080 2.910 3.550 ;
        RECT  2.470 2.060 2.710 2.800 ;
        RECT  2.390 2.560 2.470 2.800 ;
        RECT  2.150 2.560 2.390 4.340 ;
        RECT  0.830 3.010 2.150 3.250 ;
        RECT  0.500 3.010 0.830 3.380 ;
        RECT  0.570 1.390 0.810 1.830 ;
        RECT  0.500 1.590 0.570 1.830 ;
        RECT  0.430 1.590 0.500 3.380 ;
        RECT  0.260 1.590 0.430 3.250 ;
    END
END DFFRHQXL

MACRO DFFRHQX4
    CLASS CORE ;
    FOREIGN DFFRHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFRHQXL ;
    SIZE 21.120 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  14.500 1.800 14.590 2.100 ;
        RECT  14.590 1.650 15.070 2.100 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.080 2.940 18.090 3.580 ;
        RECT  18.040 0.730 18.440 1.710 ;
        RECT  18.090 2.940 18.490 3.930 ;
        RECT  18.440 1.460 19.560 1.700 ;
        RECT  18.490 2.940 19.910 3.220 ;
        RECT  19.560 0.730 19.910 1.710 ;
        RECT  19.910 0.730 19.960 3.220 ;
        RECT  19.960 1.450 20.350 3.220 ;
        RECT  20.350 2.940 20.530 3.220 ;
        RECT  20.530 2.940 20.930 3.930 ;
        RECT  20.930 2.940 20.940 3.580 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.390 2.420 1.510 3.200 ;
        RECT  1.510 2.410 1.520 3.200 ;
        RECT  1.520 2.410 1.780 3.210 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.760 1.550 1.210 2.110 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 4.480 1.390 5.440 ;
        RECT  1.390 4.640 3.520 5.440 ;
        RECT  3.520 4.480 3.920 5.440 ;
        RECT  3.920 4.640 5.280 5.440 ;
        RECT  5.280 4.480 5.680 5.440 ;
        RECT  5.680 4.640 6.940 5.440 ;
        RECT  6.940 4.070 7.180 5.440 ;
        RECT  7.180 4.640 8.480 5.440 ;
        RECT  8.480 4.480 8.880 5.440 ;
        RECT  8.880 4.640 13.770 5.440 ;
        RECT  13.770 4.190 14.010 5.440 ;
        RECT  14.010 4.640 15.330 5.440 ;
        RECT  15.330 4.480 15.730 5.440 ;
        RECT  15.730 4.640 16.940 5.440 ;
        RECT  16.940 2.840 17.360 5.440 ;
        RECT  17.360 4.640 19.310 5.440 ;
        RECT  19.310 3.730 19.710 5.440 ;
        RECT  19.710 4.640 21.120 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.010 0.400 ;
        RECT  1.010 -0.400 1.410 0.560 ;
        RECT  1.410 -0.400 3.720 0.400 ;
        RECT  3.720 -0.400 3.730 1.150 ;
        RECT  3.730 -0.400 4.130 1.350 ;
        RECT  4.130 -0.400 4.140 1.150 ;
        RECT  4.140 -0.400 5.150 0.400 ;
        RECT  5.150 -0.400 5.390 1.480 ;
        RECT  5.390 1.240 5.650 1.480 ;
        RECT  5.390 -0.400 6.760 0.400 ;
        RECT  6.760 -0.400 7.160 1.410 ;
        RECT  7.160 -0.400 8.280 0.400 ;
        RECT  8.280 -0.400 8.680 1.270 ;
        RECT  8.680 -0.400 14.080 0.400 ;
        RECT  14.080 -0.400 14.320 1.530 ;
        RECT  14.320 -0.400 15.580 0.400 ;
        RECT  15.580 -0.400 15.980 0.560 ;
        RECT  15.980 -0.400 17.360 0.400 ;
        RECT  17.360 -0.400 17.600 1.650 ;
        RECT  17.600 -0.400 18.790 0.400 ;
        RECT  18.790 -0.400 18.800 0.880 ;
        RECT  18.800 -0.400 19.200 1.080 ;
        RECT  19.200 -0.400 19.210 0.880 ;
        RECT  19.210 -0.400 20.310 0.400 ;
        RECT  20.310 -0.400 20.320 0.880 ;
        RECT  20.320 -0.400 20.720 1.080 ;
        RECT  20.720 -0.400 20.730 0.880 ;
        RECT  20.730 -0.400 21.120 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  17.080 2.120 19.470 2.360 ;
        RECT  16.840 0.860 17.080 2.570 ;
        RECT  15.080 0.860 16.840 1.100 ;
        RECT  16.670 2.170 16.840 2.570 ;
        RECT  16.580 2.170 16.670 4.180 ;
        RECT  16.430 2.250 16.580 4.180 ;
        RECT  16.320 1.380 16.560 1.780 ;
        RECT  14.910 3.940 16.430 4.180 ;
        RECT  15.630 1.540 16.320 1.780 ;
        RECT  15.910 2.170 16.150 3.660 ;
        RECT  15.050 3.420 15.910 3.660 ;
        RECT  15.390 1.540 15.630 3.140 ;
        RECT  15.330 2.370 15.390 3.140 ;
        RECT  14.010 2.370 15.330 2.610 ;
        RECT  14.840 0.860 15.080 1.360 ;
        RECT  14.810 3.150 15.050 3.660 ;
        RECT  14.530 3.940 14.910 4.230 ;
        RECT  13.490 3.150 14.810 3.390 ;
        RECT  14.510 3.670 14.530 4.230 ;
        RECT  14.290 3.670 14.510 4.180 ;
        RECT  13.490 3.670 14.290 3.910 ;
        RECT  13.770 2.210 14.010 2.610 ;
        RECT  13.370 2.210 13.770 2.450 ;
        RECT  13.250 2.730 13.490 3.390 ;
        RECT  13.250 3.670 13.490 4.370 ;
        RECT  12.980 2.730 13.250 2.970 ;
        RECT  9.400 4.130 13.250 4.370 ;
        RECT  12.740 0.670 12.980 2.970 ;
        RECT  12.730 3.250 12.970 3.850 ;
        RECT  11.550 0.670 12.740 0.910 ;
        RECT  12.370 2.570 12.740 2.970 ;
        RECT  9.920 3.610 12.730 3.850 ;
        RECT  10.730 2.570 12.370 2.810 ;
        RECT  12.140 1.190 12.300 1.430 ;
        RECT  11.900 1.190 12.140 1.810 ;
        RECT  10.450 3.090 11.950 3.330 ;
        RECT  10.780 1.570 11.900 1.810 ;
        RECT  11.540 0.670 11.550 1.210 ;
        RECT  11.140 0.670 11.540 1.330 ;
        RECT  11.130 0.670 11.140 1.210 ;
        RECT  9.560 0.670 11.130 0.910 ;
        RECT  10.450 1.190 10.780 1.810 ;
        RECT  10.210 1.190 10.450 3.330 ;
        RECT  9.360 1.190 10.210 1.430 ;
        RECT  9.910 2.820 10.210 3.140 ;
        RECT  9.690 1.740 9.930 2.440 ;
        RECT  9.680 3.420 9.920 3.850 ;
        RECT  8.740 2.820 9.910 3.060 ;
        RECT  8.220 2.200 9.690 2.440 ;
        RECT  8.220 3.420 9.680 3.660 ;
        RECT  9.160 3.940 9.400 4.370 ;
        RECT  9.120 1.190 9.360 1.790 ;
        RECT  7.700 3.940 9.160 4.180 ;
        RECT  7.840 1.550 9.120 1.790 ;
        RECT  8.500 2.740 8.740 3.140 ;
        RECT  7.980 2.200 8.220 3.660 ;
        RECT  6.920 2.200 7.980 2.440 ;
        RECT  7.600 1.110 7.840 1.790 ;
        RECT  7.460 3.390 7.700 4.180 ;
        RECT  6.400 3.390 7.460 3.630 ;
        RECT  6.680 1.770 6.920 3.110 ;
        RECT  6.320 1.770 6.680 2.010 ;
        RECT  6.370 3.910 6.610 4.310 ;
        RECT  6.160 2.290 6.400 3.630 ;
        RECT  3.310 3.940 6.370 4.180 ;
        RECT  6.080 0.670 6.320 2.010 ;
        RECT  5.570 2.290 6.160 2.530 ;
        RECT  5.670 0.670 6.080 0.910 ;
        RECT  5.290 2.930 5.880 3.330 ;
        RECT  5.050 1.770 5.290 3.330 ;
        RECT  4.870 1.770 5.050 2.010 ;
        RECT  5.030 2.950 5.050 3.330 ;
        RECT  3.830 2.950 5.030 3.190 ;
        RECT  4.630 1.070 4.870 2.010 ;
        RECT  4.350 2.290 4.670 2.530 ;
        RECT  4.570 1.070 4.630 1.470 ;
        RECT  4.110 1.750 4.350 2.530 ;
        RECT  3.280 1.750 4.110 1.990 ;
        RECT  3.590 2.270 3.830 3.190 ;
        RECT  3.040 2.580 3.310 4.180 ;
        RECT  3.040 0.920 3.280 2.300 ;
        RECT  2.360 0.920 3.040 1.160 ;
        RECT  2.590 2.060 3.040 2.300 ;
        RECT  2.870 2.580 3.040 2.980 ;
        RECT  0.570 3.940 3.040 4.180 ;
        RECT  2.590 3.260 2.710 3.660 ;
        RECT  2.350 2.060 2.590 3.660 ;
        RECT  1.800 1.500 2.430 1.740 ;
        RECT  1.560 0.860 1.800 1.740 ;
        RECT  0.590 0.860 1.560 1.100 ;
        RECT  0.490 0.670 0.590 1.100 ;
        RECT  0.490 3.040 0.570 4.180 ;
        RECT  0.250 0.670 0.490 4.180 ;
        RECT  0.190 0.670 0.250 1.070 ;
        RECT  0.170 3.040 0.250 4.180 ;
    END
END DFFRHQX4

MACRO DFFRHQX2
    CLASS CORE ;
    FOREIGN DFFRHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFRHQXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  13.310 2.730 13.750 3.220 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.310 0.990 14.710 1.390 ;
        RECT  15.160 2.960 15.380 4.050 ;
        RECT  15.380 2.950 15.510 4.050 ;
        RECT  14.710 1.150 15.510 1.390 ;
        RECT  15.510 1.150 15.560 4.050 ;
        RECT  15.560 1.150 15.640 3.210 ;
        RECT  15.640 1.150 15.750 3.200 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.210 1.290 1.450 2.350 ;
        RECT  1.450 1.290 1.520 1.530 ;
        RECT  1.520 1.270 1.780 1.530 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.740 2.660 1.130 3.210 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.980 5.440 ;
        RECT  0.980 4.480 1.380 5.440 ;
        RECT  1.380 4.640 3.320 5.440 ;
        RECT  3.320 4.310 3.330 5.440 ;
        RECT  3.330 4.190 3.730 5.440 ;
        RECT  3.730 4.310 3.740 5.440 ;
        RECT  3.740 4.640 7.230 5.440 ;
        RECT  7.230 4.480 7.630 5.440 ;
        RECT  7.630 4.640 10.950 5.440 ;
        RECT  10.950 4.480 11.350 5.440 ;
        RECT  12.760 3.180 13.000 3.730 ;
        RECT  11.350 4.640 14.020 5.440 ;
        RECT  13.000 3.490 14.020 3.730 ;
        RECT  14.020 3.490 14.260 5.440 ;
        RECT  14.260 4.640 16.370 5.440 ;
        RECT  16.370 3.650 16.380 5.440 ;
        RECT  16.380 3.160 16.780 5.440 ;
        RECT  16.780 3.650 16.790 5.440 ;
        RECT  16.790 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.030 0.400 ;
        RECT  1.030 -0.400 1.430 0.560 ;
        RECT  1.430 -0.400 3.360 0.400 ;
        RECT  3.360 -0.400 3.520 1.170 ;
        RECT  3.520 -0.400 3.760 1.440 ;
        RECT  3.760 1.200 4.910 1.440 ;
        RECT  4.910 1.200 5.310 1.600 ;
        RECT  3.760 -0.400 7.380 0.400 ;
        RECT  7.380 -0.400 7.390 0.940 ;
        RECT  7.390 -0.400 7.790 1.060 ;
        RECT  7.790 -0.400 7.800 0.940 ;
        RECT  7.800 -0.400 11.320 0.400 ;
        RECT  11.320 -0.400 11.720 0.560 ;
        RECT  11.720 -0.400 12.900 0.400 ;
        RECT  12.900 -0.400 13.880 0.560 ;
        RECT  13.880 -0.400 15.060 0.400 ;
        RECT  15.060 -0.400 15.070 0.750 ;
        RECT  15.070 -0.400 15.470 0.870 ;
        RECT  15.470 -0.400 15.480 0.750 ;
        RECT  15.480 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  15.070 1.990 15.230 2.390 ;
        RECT  14.830 1.670 15.070 2.390 ;
        RECT  14.030 1.670 14.830 1.910 ;
        RECT  13.280 2.200 14.460 2.440 ;
        RECT  13.790 0.860 14.030 1.910 ;
        RECT  12.070 0.860 13.790 1.100 ;
        RECT  12.400 4.050 13.580 4.290 ;
        RECT  12.880 1.630 13.280 2.440 ;
        RECT  12.840 2.200 12.880 2.440 ;
        RECT  12.520 2.200 12.840 2.660 ;
        RECT  12.400 2.420 12.520 2.660 ;
        RECT  11.700 1.470 12.420 1.710 ;
        RECT  12.160 2.420 12.400 4.290 ;
        RECT  10.290 3.940 12.160 4.180 ;
        RECT  11.670 0.860 12.070 1.150 ;
        RECT  11.700 3.160 11.860 3.400 ;
        RECT  11.460 1.470 11.700 3.400 ;
        RECT  10.380 0.860 11.670 1.100 ;
        RECT  11.180 2.590 11.460 2.830 ;
        RECT  10.380 1.480 10.620 2.900 ;
        RECT  9.980 0.710 10.380 1.100 ;
        RECT  10.280 2.660 10.380 2.900 ;
        RECT  10.050 3.940 10.290 4.370 ;
        RECT  10.040 2.660 10.280 3.060 ;
        RECT  9.810 1.450 10.050 2.380 ;
        RECT  8.150 4.130 10.050 4.370 ;
        RECT  9.770 3.390 10.030 3.630 ;
        RECT  9.290 0.860 9.980 1.100 ;
        RECT  9.710 2.140 9.810 2.380 ;
        RECT  9.710 3.390 9.770 3.850 ;
        RECT  9.470 2.140 9.710 3.850 ;
        RECT  8.670 3.610 9.470 3.850 ;
        RECT  9.190 0.860 9.290 1.850 ;
        RECT  9.050 0.860 9.190 3.330 ;
        RECT  8.950 1.610 9.050 3.330 ;
        RECT  8.610 1.340 8.670 3.850 ;
        RECT  8.430 1.150 8.610 3.850 ;
        RECT  8.210 1.150 8.430 1.580 ;
        RECT  6.750 3.420 8.430 3.660 ;
        RECT  7.110 1.340 8.210 1.580 ;
        RECT  7.910 2.150 8.150 2.550 ;
        RECT  7.910 3.940 8.150 4.370 ;
        RECT  7.130 2.230 7.910 2.470 ;
        RECT  5.450 3.940 7.910 4.180 ;
        RECT  6.890 1.860 7.130 3.140 ;
        RECT  6.870 1.040 7.110 1.580 ;
        RECT  6.490 1.860 6.890 2.100 ;
        RECT  6.410 2.900 6.890 3.140 ;
        RECT  6.570 1.040 6.870 1.280 ;
        RECT  5.970 2.380 6.610 2.620 ;
        RECT  6.290 1.560 6.490 2.100 ;
        RECT  6.170 2.900 6.410 3.430 ;
        RECT  6.250 1.200 6.290 2.100 ;
        RECT  6.050 1.200 6.250 1.800 ;
        RECT  6.010 3.190 6.170 3.430 ;
        RECT  5.810 0.680 6.050 1.440 ;
        RECT  5.730 2.080 5.970 2.620 ;
        RECT  4.050 0.680 5.810 0.920 ;
        RECT  4.690 2.080 5.730 2.320 ;
        RECT  5.210 2.600 5.450 4.180 ;
        RECT  5.050 2.600 5.210 2.840 ;
        RECT  4.450 2.080 4.690 3.590 ;
        RECT  4.440 2.080 4.450 2.320 ;
        RECT  4.410 3.350 4.450 3.590 ;
        RECT  4.430 1.840 4.440 2.320 ;
        RECT  4.030 1.720 4.430 2.320 ;
        RECT  4.170 3.350 4.410 3.750 ;
        RECT  4.090 2.600 4.170 2.840 ;
        RECT  3.770 2.600 4.090 3.060 ;
        RECT  4.020 1.840 4.030 2.320 ;
        RECT  3.330 2.080 4.020 2.320 ;
        RECT  2.790 2.820 3.770 3.060 ;
        RECT  3.090 2.080 3.330 2.540 ;
        RECT  2.530 3.940 2.930 4.210 ;
        RECT  2.750 2.820 2.790 3.520 ;
        RECT  2.510 0.670 2.750 3.520 ;
        RECT  2.030 3.940 2.530 4.180 ;
        RECT  1.990 0.670 2.510 0.910 ;
        RECT  2.310 3.120 2.510 3.520 ;
        RECT  2.030 1.940 2.170 2.840 ;
        RECT  1.930 1.940 2.030 4.180 ;
        RECT  1.790 2.600 1.930 4.180 ;
        RECT  0.570 3.490 1.790 3.730 ;
        RECT  0.410 1.370 0.570 1.770 ;
        RECT  0.410 3.490 0.570 3.890 ;
        RECT  0.170 1.370 0.410 3.890 ;
    END
END DFFRHQX2

MACRO DFFRHQX1
    CLASS CORE ;
    FOREIGN DFFRHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFRHQXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  11.770 2.910 12.430 3.260 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.480 0.780 12.650 1.020 ;
        RECT  12.650 0.780 12.890 1.480 ;
        RECT  13.350 2.950 13.460 3.830 ;
        RECT  12.890 1.240 13.460 1.480 ;
        RECT  13.460 1.240 13.700 3.830 ;
        RECT  13.700 2.950 13.710 3.830 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 1.700 1.500 2.100 ;
        RECT  1.500 1.700 1.620 2.200 ;
        RECT  1.620 1.700 1.870 2.210 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.770 2.380 1.120 2.930 ;
        RECT  1.120 2.520 1.300 2.920 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.530 5.440 ;
        RECT  1.530 3.940 1.770 5.440 ;
        RECT  1.770 4.640 3.660 5.440 ;
        RECT  3.660 4.140 3.670 5.440 ;
        RECT  3.670 4.020 4.070 5.440 ;
        RECT  4.070 4.140 4.080 5.440 ;
        RECT  4.080 4.640 6.890 5.440 ;
        RECT  6.890 4.480 7.290 5.440 ;
        RECT  7.290 4.640 9.810 5.440 ;
        RECT  9.810 4.480 10.210 5.440 ;
        RECT  11.100 3.070 11.260 3.310 ;
        RECT  11.260 3.070 11.500 3.770 ;
        RECT  10.210 4.640 12.140 5.440 ;
        RECT  11.500 3.530 12.140 3.770 ;
        RECT  12.140 3.530 12.380 5.440 ;
        RECT  12.380 4.640 13.860 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.320 0.400 ;
        RECT  1.320 -0.400 1.720 0.560 ;
        RECT  1.720 -0.400 3.620 0.400 ;
        RECT  3.620 -0.400 3.630 0.860 ;
        RECT  3.630 -0.400 3.790 0.980 ;
        RECT  3.790 -0.400 4.030 1.440 ;
        RECT  4.030 -0.400 4.040 0.860 ;
        RECT  4.030 1.200 5.170 1.440 ;
        RECT  5.170 1.200 5.410 1.760 ;
        RECT  5.410 1.520 5.650 1.760 ;
        RECT  4.040 -0.400 6.650 0.400 ;
        RECT  6.650 -0.400 6.890 1.160 ;
        RECT  6.890 -0.400 9.500 0.400 ;
        RECT  9.500 -0.400 9.900 0.560 ;
        RECT  9.900 -0.400 11.140 0.400 ;
        RECT  11.140 -0.400 11.540 0.560 ;
        RECT  11.540 -0.400 13.270 0.400 ;
        RECT  13.270 -0.400 13.280 0.760 ;
        RECT  13.280 -0.400 13.680 0.960 ;
        RECT  13.680 -0.400 13.690 0.760 ;
        RECT  13.690 -0.400 13.860 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.020 1.760 13.180 2.000 ;
        RECT  12.700 2.400 12.940 2.810 ;
        RECT  11.300 2.400 12.700 2.640 ;
        RECT  11.780 0.860 12.020 2.000 ;
        RECT  10.410 0.860 11.780 1.100 ;
        RECT  10.740 4.050 11.700 4.290 ;
        RECT  11.300 1.380 11.460 1.620 ;
        RECT  11.060 1.380 11.300 2.640 ;
        RECT  10.740 2.130 11.060 2.370 ;
        RECT  10.500 2.130 10.740 4.290 ;
        RECT  10.060 1.470 10.610 1.710 ;
        RECT  5.790 3.940 10.500 4.180 ;
        RECT  9.860 0.860 10.410 1.150 ;
        RECT  10.060 3.210 10.220 3.450 ;
        RECT  9.820 1.470 10.060 3.450 ;
        RECT  9.400 0.860 9.860 1.100 ;
        RECT  9.700 2.550 9.820 2.950 ;
        RECT  9.160 0.860 9.400 2.350 ;
        RECT  8.470 0.860 9.160 1.110 ;
        RECT  9.150 2.110 9.160 2.350 ;
        RECT  8.910 2.110 9.150 3.660 ;
        RECT  8.470 3.420 8.910 3.660 ;
        RECT  8.630 1.590 8.880 1.830 ;
        RECT  8.390 1.590 8.630 3.140 ;
        RECT  8.230 0.860 8.470 1.310 ;
        RECT  7.910 1.590 8.110 3.660 ;
        RECT  7.870 1.060 7.910 3.660 ;
        RECT  7.670 1.060 7.870 1.830 ;
        RECT  7.710 3.420 7.870 3.660 ;
        RECT  7.390 1.060 7.670 1.300 ;
        RECT  7.390 2.300 7.590 2.700 ;
        RECT  7.150 1.580 7.390 3.660 ;
        RECT  6.170 1.580 7.150 1.820 ;
        RECT  6.410 3.420 7.150 3.660 ;
        RECT  6.630 2.170 6.870 3.140 ;
        RECT  4.890 2.170 6.630 2.410 ;
        RECT  5.930 0.680 6.170 1.820 ;
        RECT  4.310 0.680 5.930 0.920 ;
        RECT  5.550 2.690 5.790 4.180 ;
        RECT  5.390 2.690 5.550 2.930 ;
        RECT  4.650 1.720 4.890 3.710 ;
        RECT  3.650 1.720 4.650 1.960 ;
        RECT  4.510 3.310 4.650 3.710 ;
        RECT  4.130 2.550 4.370 2.950 ;
        RECT  2.980 2.710 4.130 2.950 ;
        RECT  3.410 1.720 3.650 2.400 ;
        RECT  2.370 3.820 3.270 4.060 ;
        RECT  2.740 0.670 2.980 3.540 ;
        RECT  2.290 0.670 2.740 0.910 ;
        RECT  2.650 3.140 2.740 3.540 ;
        RECT  2.370 1.800 2.460 2.860 ;
        RECT  2.220 1.800 2.370 4.060 ;
        RECT  2.130 2.620 2.220 4.060 ;
        RECT  0.500 3.200 2.130 3.440 ;
        RECT  0.500 1.220 0.860 1.620 ;
        RECT  0.460 1.220 0.500 3.440 ;
        RECT  0.260 1.380 0.460 3.440 ;
    END
END DFFRHQX1

MACRO DFFRXL
    CLASS CORE ;
    FOREIGN DFFRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.520 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.060 2.850 4.590 3.260 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.600 3.670 12.740 4.070 ;
        RECT  12.740 3.510 13.080 4.070 ;
        RECT  12.690 0.730 13.090 1.100 ;
        RECT  13.080 3.520 13.430 3.760 ;
        RECT  13.090 0.860 13.430 1.100 ;
        RECT  13.430 0.860 13.670 3.760 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.950 1.390 13.970 1.790 ;
        RECT  13.970 1.390 14.060 1.820 ;
        RECT  13.950 2.980 14.070 3.380 ;
        RECT  14.060 1.390 14.070 2.090 ;
        RECT  14.070 1.390 14.190 3.380 ;
        RECT  14.190 1.500 14.300 3.380 ;
        RECT  14.300 1.830 14.310 3.380 ;
        RECT  14.310 1.830 14.320 2.090 ;
        RECT  14.310 2.980 14.350 3.380 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.950 1.590 3.210 ;
        RECT  1.590 2.530 1.780 3.210 ;
        RECT  1.780 2.530 1.830 3.200 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.480 2.270 0.880 2.670 ;
        RECT  0.880 2.390 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.080 5.440 ;
        RECT  1.080 4.480 1.480 5.440 ;
        RECT  1.480 4.640 3.430 5.440 ;
        RECT  3.430 4.480 3.830 5.440 ;
        RECT  3.830 4.640 7.000 5.440 ;
        RECT  7.000 4.110 7.980 5.440 ;
        RECT  7.980 4.640 9.850 5.440 ;
        RECT  9.850 4.170 9.860 5.440 ;
        RECT  9.860 3.970 10.260 5.440 ;
        RECT  10.260 4.170 10.270 5.440 ;
        RECT  10.270 4.640 11.830 5.440 ;
        RECT  11.830 3.860 11.840 5.440 ;
        RECT  11.840 3.660 12.240 5.440 ;
        RECT  12.240 3.860 12.250 5.440 ;
        RECT  12.250 4.640 13.340 5.440 ;
        RECT  13.340 4.480 13.740 5.440 ;
        RECT  13.740 4.640 14.520 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        RECT  0.940 -0.400 1.340 0.560 ;
        RECT  1.340 -0.400 3.540 0.400 ;
        RECT  3.540 -0.400 3.550 0.730 ;
        RECT  3.550 -0.400 3.950 0.850 ;
        RECT  3.950 -0.400 3.960 0.730 ;
        RECT  3.960 -0.400 5.570 0.400 ;
        RECT  5.570 -0.400 5.830 1.530 ;
        RECT  5.830 1.290 7.350 1.530 ;
        RECT  7.350 1.290 7.590 1.840 ;
        RECT  7.590 1.440 7.750 1.840 ;
        RECT  5.830 -0.400 10.040 0.400 ;
        RECT  10.040 -0.400 10.440 1.290 ;
        RECT  10.440 -0.400 11.790 0.400 ;
        RECT  11.790 -0.400 11.800 0.890 ;
        RECT  11.800 -0.400 12.200 1.090 ;
        RECT  12.200 -0.400 12.210 0.890 ;
        RECT  12.210 -0.400 13.750 0.400 ;
        RECT  13.750 -0.400 14.150 0.560 ;
        RECT  14.150 -0.400 14.520 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.910 1.470 13.150 3.150 ;
        RECT  12.690 1.470 12.910 1.710 ;
        RECT  12.610 2.750 12.910 3.150 ;
        RECT  11.680 1.970 12.360 2.370 ;
        RECT  11.440 1.590 11.680 3.270 ;
        RECT  11.320 1.590 11.440 1.830 ;
        RECT  11.020 3.030 11.440 3.270 ;
        RECT  10.920 0.890 11.320 1.830 ;
        RECT  10.760 2.110 11.160 2.510 ;
        RECT  10.780 3.030 11.020 4.010 ;
        RECT  10.160 1.590 10.920 1.830 ;
        RECT  10.620 3.610 10.780 4.010 ;
        RECT  9.480 2.270 10.760 2.510 ;
        RECT  9.760 1.590 10.160 1.990 ;
        RECT  9.480 3.730 9.520 4.130 ;
        RECT  9.470 2.270 9.480 4.130 ;
        RECT  9.230 1.180 9.470 4.130 ;
        RECT  9.100 1.180 9.230 1.420 ;
        RECT  9.120 3.730 9.230 4.130 ;
        RECT  8.700 1.020 9.100 1.420 ;
        RECT  8.840 2.380 8.920 2.780 ;
        RECT  8.600 2.380 8.840 3.830 ;
        RECT  8.320 1.740 8.800 1.980 ;
        RECT  7.120 3.590 8.600 3.830 ;
        RECT  8.080 0.670 8.320 3.310 ;
        RECT  6.110 0.670 8.080 0.910 ;
        RECT  7.400 3.070 8.080 3.310 ;
        RECT  6.470 2.160 7.800 2.560 ;
        RECT  6.880 2.880 7.120 3.830 ;
        RECT  6.410 3.590 6.880 3.830 ;
        RECT  6.230 1.820 6.470 3.140 ;
        RECT  6.170 3.590 6.410 4.290 ;
        RECT  5.290 1.820 6.230 2.060 ;
        RECT  5.780 2.900 6.230 3.140 ;
        RECT  4.360 4.050 6.170 4.290 ;
        RECT  5.100 2.340 5.950 2.580 ;
        RECT  5.540 2.900 5.780 3.770 ;
        RECT  5.380 3.530 5.540 3.770 ;
        RECT  5.160 1.650 5.290 2.060 ;
        RECT  5.050 1.120 5.160 2.060 ;
        RECT  4.860 2.340 5.100 3.770 ;
        RECT  4.920 1.120 5.050 1.890 ;
        RECT  3.650 1.650 4.920 1.890 ;
        RECT  4.770 2.340 4.860 2.580 ;
        RECT  4.640 3.530 4.860 3.770 ;
        RECT  4.370 2.170 4.770 2.580 ;
        RECT  4.470 0.770 4.640 1.010 ;
        RECT  4.230 0.770 4.470 1.370 ;
        RECT  4.120 3.940 4.360 4.290 ;
        RECT  2.910 1.130 4.230 1.370 ;
        RECT  3.150 3.940 4.120 4.180 ;
        RECT  3.410 1.650 3.650 2.830 ;
        RECT  3.250 2.430 3.410 2.830 ;
        RECT  2.750 3.940 3.150 4.370 ;
        RECT  2.670 1.130 2.910 3.650 ;
        RECT  2.390 3.940 2.750 4.180 ;
        RECT  2.210 1.130 2.670 1.550 ;
        RECT  2.150 1.890 2.390 4.180 ;
        RECT  1.910 1.890 2.150 2.130 ;
        RECT  2.100 3.510 2.150 4.180 ;
        RECT  0.570 3.510 2.100 3.750 ;
        RECT  1.670 1.410 1.910 2.130 ;
        RECT  0.570 1.410 1.670 1.650 ;
        RECT  0.170 1.250 0.570 1.650 ;
        RECT  0.170 3.350 0.570 3.750 ;
    END
END DFFRXL

MACRO DFFRX4
    CLASS CORE ;
    FOREIGN DFFRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFRXL ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.010 2.610 4.020 3.050 ;
        RECT  4.020 2.610 4.420 3.210 ;
        RECT  4.420 2.610 4.430 3.050 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.040 2.750 17.270 3.150 ;
        RECT  17.030 1.170 17.270 1.570 ;
        RECT  17.270 1.170 17.670 3.220 ;
        RECT  17.670 1.820 17.710 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.580 2.750 18.590 3.150 ;
        RECT  18.570 1.170 18.590 1.570 ;
        RECT  18.590 1.170 18.970 3.150 ;
        RECT  18.970 1.260 18.990 3.150 ;
        RECT  18.990 1.260 19.030 2.660 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.250 1.300 1.490 2.090 ;
        RECT  1.490 1.300 1.520 1.540 ;
        RECT  1.520 1.270 1.770 1.540 ;
        RECT  1.770 1.270 1.780 1.530 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.770 2.500 0.780 2.920 ;
        RECT  0.780 2.400 0.860 2.920 ;
        RECT  0.860 2.390 1.120 2.920 ;
        RECT  1.120 2.500 1.190 2.920 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.910 5.440 ;
        RECT  0.910 4.480 1.310 5.440 ;
        RECT  1.310 4.640 3.590 5.440 ;
        RECT  3.590 4.480 3.990 5.440 ;
        RECT  3.990 4.640 7.170 5.440 ;
        RECT  7.170 4.180 8.710 5.440 ;
        RECT  8.710 4.640 11.250 5.440 ;
        RECT  11.250 4.290 11.260 5.440 ;
        RECT  11.260 4.090 11.660 5.440 ;
        RECT  11.660 4.290 11.670 5.440 ;
        RECT  11.670 4.640 12.580 5.440 ;
        RECT  12.580 4.080 12.980 5.440 ;
        RECT  12.980 4.640 15.010 5.440 ;
        RECT  15.010 2.960 15.410 5.440 ;
        RECT  15.410 4.640 16.350 5.440 ;
        RECT  16.350 4.480 16.750 5.440 ;
        RECT  16.750 4.640 17.860 5.440 ;
        RECT  17.860 4.210 17.870 5.440 ;
        RECT  17.870 4.010 18.270 5.440 ;
        RECT  18.270 4.210 18.280 5.440 ;
        RECT  18.280 4.640 19.220 5.440 ;
        RECT  19.220 4.210 19.230 5.440 ;
        RECT  19.230 4.010 19.630 5.440 ;
        RECT  19.630 4.210 19.640 5.440 ;
        RECT  19.640 4.640 19.800 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.040 0.400 ;
        RECT  1.040 -0.400 1.440 0.560 ;
        RECT  1.440 -0.400 4.370 0.400 ;
        RECT  4.370 -0.400 5.350 1.290 ;
        RECT  5.350 -0.400 6.280 0.400 ;
        RECT  6.280 -0.400 6.290 0.890 ;
        RECT  6.290 -0.400 6.690 1.090 ;
        RECT  6.690 -0.400 6.700 0.890 ;
        RECT  6.700 -0.400 7.990 0.400 ;
        RECT  7.990 -0.400 8.000 1.120 ;
        RECT  8.000 -0.400 8.400 1.320 ;
        RECT  8.400 -0.400 8.410 1.120 ;
        RECT  8.410 -0.400 10.580 0.400 ;
        RECT  10.580 -0.400 10.980 1.090 ;
        RECT  10.980 -0.400 12.880 0.400 ;
        RECT  12.880 -0.400 13.860 1.010 ;
        RECT  13.860 -0.400 14.910 0.400 ;
        RECT  14.910 -0.400 15.310 1.620 ;
        RECT  15.310 -0.400 16.420 0.400 ;
        RECT  16.420 -0.400 16.820 0.890 ;
        RECT  16.820 -0.400 17.850 0.400 ;
        RECT  17.850 -0.400 17.860 0.690 ;
        RECT  17.860 -0.400 18.260 0.890 ;
        RECT  18.260 -0.400 18.270 0.690 ;
        RECT  18.270 -0.400 19.210 0.400 ;
        RECT  19.210 -0.400 19.220 0.690 ;
        RECT  19.220 -0.400 19.620 0.890 ;
        RECT  19.620 -0.400 19.630 0.690 ;
        RECT  19.630 -0.400 19.800 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  19.270 2.180 19.510 3.730 ;
        RECT  16.630 3.490 19.270 3.730 ;
        RECT  16.390 1.550 16.630 3.730 ;
        RECT  16.100 1.550 16.390 1.790 ;
        RECT  15.730 3.330 16.390 3.730 ;
        RECT  14.590 2.070 16.150 2.470 ;
        RECT  15.700 1.390 16.100 1.790 ;
        RECT  14.350 0.660 14.590 3.490 ;
        RECT  14.190 0.660 14.350 1.640 ;
        RECT  14.230 3.250 14.350 3.490 ;
        RECT  14.150 3.250 14.230 3.650 ;
        RECT  12.880 1.390 14.190 1.630 ;
        RECT  13.830 3.250 14.150 3.790 ;
        RECT  13.710 2.200 14.110 2.600 ;
        RECT  12.300 3.550 13.830 3.790 ;
        RECT  12.400 2.200 13.710 2.530 ;
        RECT  12.640 1.250 12.880 1.630 ;
        RECT  12.480 1.250 12.640 1.490 ;
        RECT  12.240 2.130 12.400 2.530 ;
        RECT  12.060 3.550 12.300 4.350 ;
        RECT  12.000 1.650 12.240 3.270 ;
        RECT  11.800 1.650 12.000 1.890 ;
        RECT  11.610 3.030 12.000 3.270 ;
        RECT  11.560 0.680 11.800 1.890 ;
        RECT  11.480 2.340 11.720 2.740 ;
        RECT  11.370 3.030 11.610 3.450 ;
        RECT  11.330 0.680 11.560 1.620 ;
        RECT  11.280 2.340 11.480 2.580 ;
        RECT  10.380 3.210 11.370 3.450 ;
        RECT  10.100 1.380 11.330 1.620 ;
        RECT  11.040 1.900 11.280 2.580 ;
        RECT  9.380 1.900 11.040 2.140 ;
        RECT  9.590 2.690 10.630 2.930 ;
        RECT  10.140 3.210 10.380 3.860 ;
        RECT  9.980 3.460 10.140 3.860 ;
        RECT  9.860 1.190 10.100 1.620 ;
        RECT  9.220 1.190 9.860 1.430 ;
        RECT  9.350 2.690 9.590 3.900 ;
        RECT  9.300 1.730 9.380 2.140 ;
        RECT  7.710 3.660 9.350 3.900 ;
        RECT  9.060 1.710 9.300 2.140 ;
        RECT  8.820 1.710 9.060 3.160 ;
        RECT  7.440 1.710 8.820 1.950 ;
        RECT  8.230 2.920 8.820 3.160 ;
        RECT  6.880 2.250 8.540 2.490 ;
        RECT  7.990 2.920 8.230 3.380 ;
        RECT  7.470 2.770 7.710 3.900 ;
        RECT  7.310 2.770 7.470 3.540 ;
        RECT  7.200 0.670 7.440 1.950 ;
        RECT  6.810 3.300 7.310 3.540 ;
        RECT  6.980 0.670 7.200 0.910 ;
        RECT  6.640 1.570 6.880 3.020 ;
        RECT  6.570 3.300 6.810 4.270 ;
        RECT  3.540 1.570 6.640 1.810 ;
        RECT  6.290 2.780 6.640 3.020 ;
        RECT  4.510 4.030 6.570 4.270 ;
        RECT  5.030 2.150 6.360 2.390 ;
        RECT  6.050 2.780 6.290 3.690 ;
        RECT  5.890 3.450 6.050 3.690 ;
        RECT  5.030 3.510 5.360 3.750 ;
        RECT  4.790 2.090 5.030 3.750 ;
        RECT  4.780 2.090 4.790 2.390 ;
        RECT  4.340 2.090 4.780 2.330 ;
        RECT  4.270 3.940 4.510 4.270 ;
        RECT  3.310 3.940 4.270 4.180 ;
        RECT  2.860 0.770 4.100 1.010 ;
        RECT  3.540 2.290 3.550 2.690 ;
        RECT  3.310 1.570 3.540 2.690 ;
        RECT  3.300 1.570 3.310 2.530 ;
        RECT  3.070 3.940 3.310 4.350 ;
        RECT  1.990 4.110 3.070 4.350 ;
        RECT  2.620 0.770 2.860 3.660 ;
        RECT  2.180 1.110 2.620 1.510 ;
        RECT  2.510 3.420 2.620 3.660 ;
        RECT  2.270 3.420 2.510 3.830 ;
        RECT  1.990 1.880 2.180 3.050 ;
        RECT  1.940 1.880 1.990 4.350 ;
        RECT  1.750 2.810 1.940 4.350 ;
        RECT  0.620 3.420 1.750 3.660 ;
        RECT  0.460 3.330 0.620 3.730 ;
        RECT  0.460 1.100 0.580 1.500 ;
        RECT  0.220 1.100 0.460 3.730 ;
        RECT  0.180 1.100 0.220 1.500 ;
    END
END DFFRX4

MACRO DFFRX2
    CLASS CORE ;
    FOREIGN DFFRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFRXL ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 2.950 3.510 3.210 ;
        RECT  3.510 2.710 3.760 3.210 ;
        RECT  3.760 2.710 4.260 3.110 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.740 2.920 13.820 3.320 ;
        RECT  13.820 2.610 13.830 3.320 ;
        RECT  13.740 0.730 13.830 1.710 ;
        RECT  13.830 0.730 14.070 3.320 ;
        RECT  14.070 2.390 14.140 3.320 ;
        RECT  14.070 0.730 14.140 1.710 ;
        RECT  14.140 2.390 14.320 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.270 0.730 15.290 1.710 ;
        RECT  15.290 0.730 15.380 1.820 ;
        RECT  15.270 3.170 15.390 4.150 ;
        RECT  15.380 0.730 15.390 2.090 ;
        RECT  15.390 0.730 15.630 4.150 ;
        RECT  15.630 0.730 15.640 2.090 ;
        RECT  15.630 3.170 15.670 4.150 ;
        RECT  15.640 0.730 15.670 1.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.380 1.150 2.660 ;
        RECT  1.150 2.320 1.490 2.740 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.510 2.420 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.870 5.440 ;
        RECT  0.870 4.480 1.270 5.440 ;
        RECT  1.270 4.640 3.350 5.440 ;
        RECT  3.350 4.480 3.750 5.440 ;
        RECT  3.750 4.640 6.650 5.440 ;
        RECT  6.650 4.170 8.190 5.440 ;
        RECT  8.190 4.640 10.210 5.440 ;
        RECT  10.210 4.110 10.220 5.440 ;
        RECT  10.220 3.910 10.620 5.440 ;
        RECT  10.620 4.110 10.630 5.440 ;
        RECT  10.630 4.640 12.170 5.440 ;
        RECT  12.170 3.500 12.180 5.440 ;
        RECT  12.180 3.300 12.580 5.440 ;
        RECT  12.580 3.500 12.590 5.440 ;
        RECT  12.590 4.640 14.500 5.440 ;
        RECT  14.500 4.320 14.510 5.440 ;
        RECT  14.510 4.120 14.910 5.440 ;
        RECT  14.910 4.320 14.920 5.440 ;
        RECT  14.920 4.640 15.840 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.740 0.400 ;
        RECT  0.740 -0.400 1.140 0.560 ;
        RECT  1.140 -0.400 4.210 0.400 ;
        RECT  4.210 -0.400 4.610 1.310 ;
        RECT  4.610 -0.400 5.700 0.400 ;
        RECT  5.700 -0.400 5.710 0.640 ;
        RECT  5.710 -0.400 6.110 0.930 ;
        RECT  6.110 -0.400 6.120 0.640 ;
        RECT  6.120 -0.400 7.400 0.400 ;
        RECT  7.400 -0.400 7.410 1.020 ;
        RECT  7.410 -0.400 7.810 1.140 ;
        RECT  7.810 -0.400 7.820 1.020 ;
        RECT  7.820 -0.400 10.490 0.400 ;
        RECT  10.490 -0.400 10.890 0.560 ;
        RECT  10.890 -0.400 12.060 0.400 ;
        RECT  12.060 -0.400 12.070 1.100 ;
        RECT  12.070 -0.400 12.470 1.300 ;
        RECT  12.470 -0.400 12.480 1.100 ;
        RECT  12.480 -0.400 14.500 0.400 ;
        RECT  14.500 -0.400 14.510 1.200 ;
        RECT  14.510 -0.400 14.910 1.690 ;
        RECT  14.910 -0.400 14.920 1.200 ;
        RECT  14.920 -0.400 15.840 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.990 2.200 15.020 2.600 ;
        RECT  14.750 2.200 14.990 3.840 ;
        RECT  13.460 3.600 14.750 3.840 ;
        RECT  13.220 1.080 13.460 3.840 ;
        RECT  12.890 1.080 13.220 1.480 ;
        RECT  13.000 2.920 13.220 3.320 ;
        RECT  11.990 1.950 12.980 2.350 ;
        RECT  11.750 1.580 11.990 3.020 ;
        RECT  11.710 1.580 11.750 1.820 ;
        RECT  11.360 2.780 11.750 3.020 ;
        RECT  11.310 0.940 11.710 1.820 ;
        RECT  11.070 2.100 11.470 2.500 ;
        RECT  11.120 2.780 11.360 3.900 ;
        RECT  10.440 1.580 11.310 1.820 ;
        RECT  10.960 2.920 11.120 3.900 ;
        RECT  9.760 2.260 11.070 2.500 ;
        RECT  10.040 1.580 10.440 1.980 ;
        RECT  9.520 1.260 9.760 3.490 ;
        RECT  9.090 1.260 9.520 1.500 ;
        RECT  9.400 3.250 9.520 3.490 ;
        RECT  9.160 3.250 9.400 3.650 ;
        RECT  8.820 2.610 9.240 2.850 ;
        RECT  8.690 1.100 9.090 1.500 ;
        RECT  8.300 1.890 8.830 2.130 ;
        RECT  8.580 2.610 8.820 3.890 ;
        RECT  6.960 3.650 8.580 3.890 ;
        RECT  8.060 1.420 8.300 3.350 ;
        RECT  6.930 1.420 8.060 1.710 ;
        RECT  7.240 3.110 8.060 3.350 ;
        RECT  7.580 1.990 7.820 2.710 ;
        RECT  6.190 1.990 7.580 2.230 ;
        RECT  6.960 2.510 7.140 2.750 ;
        RECT  6.720 2.510 6.960 3.890 ;
        RECT  6.800 1.310 6.930 1.710 ;
        RECT  6.790 0.880 6.800 1.710 ;
        RECT  6.530 0.670 6.790 1.710 ;
        RECT  6.280 3.650 6.720 3.890 ;
        RECT  6.390 0.670 6.530 0.910 ;
        RECT  6.040 3.650 6.280 4.310 ;
        RECT  5.950 1.590 6.190 3.190 ;
        RECT  4.270 4.070 6.040 4.310 ;
        RECT  5.530 1.590 5.950 1.830 ;
        RECT  5.720 2.950 5.950 3.190 ;
        RECT  5.480 2.950 5.720 3.790 ;
        RECT  5.430 2.110 5.670 2.510 ;
        RECT  5.130 1.270 5.530 1.830 ;
        RECT  5.320 3.390 5.480 3.790 ;
        RECT  4.790 2.110 5.430 2.350 ;
        RECT  3.480 1.590 5.130 1.830 ;
        RECT  4.550 2.110 4.790 3.790 ;
        RECT  4.250 2.110 4.550 2.350 ;
        RECT  4.030 3.940 4.270 4.310 ;
        RECT  3.050 3.940 4.030 4.180 ;
        RECT  3.690 0.690 3.930 1.090 ;
        RECT  2.800 0.850 3.690 1.090 ;
        RECT  3.240 1.590 3.480 2.280 ;
        RECT  3.080 1.880 3.240 2.280 ;
        RECT  2.810 3.940 3.050 4.250 ;
        RECT  2.010 4.010 2.810 4.250 ;
        RECT  2.560 0.850 2.800 3.330 ;
        RECT  2.460 0.850 2.560 1.090 ;
        RECT  2.530 3.090 2.560 3.330 ;
        RECT  2.290 3.090 2.530 3.490 ;
        RECT  2.060 0.750 2.460 1.090 ;
        RECT  2.010 1.800 2.200 2.290 ;
        RECT  1.770 1.800 2.010 4.250 ;
        RECT  1.720 1.800 1.770 2.040 ;
        RECT  0.170 3.490 1.770 3.730 ;
        RECT  1.480 1.310 1.720 2.040 ;
        RECT  0.170 1.310 1.480 1.550 ;
    END
END DFFRX2

MACRO DFFRX1
    CLASS CORE ;
    FOREIGN DFFRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFRXL ;
    SIZE 14.520 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.060 2.850 4.590 3.260 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.600 3.670 12.740 4.070 ;
        RECT  12.540 0.710 12.950 1.100 ;
        RECT  12.740 3.510 13.080 4.070 ;
        RECT  13.080 3.520 13.430 3.760 ;
        RECT  12.950 0.860 13.430 1.100 ;
        RECT  13.430 0.860 13.670 3.760 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.950 1.320 13.970 1.720 ;
        RECT  13.970 1.320 14.060 1.820 ;
        RECT  13.950 2.980 14.070 3.380 ;
        RECT  14.060 1.320 14.070 2.090 ;
        RECT  14.070 1.320 14.310 3.380 ;
        RECT  14.310 1.320 14.320 2.090 ;
        RECT  14.310 2.980 14.350 3.380 ;
        RECT  14.320 1.320 14.350 1.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.500 1.870 3.220 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.750 2.380 1.120 2.890 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.130 5.440 ;
        RECT  1.130 4.480 1.530 5.440 ;
        RECT  1.530 4.640 3.430 5.440 ;
        RECT  3.430 4.480 3.830 5.440 ;
        RECT  3.830 4.640 7.000 5.440 ;
        RECT  7.000 4.110 7.980 5.440 ;
        RECT  7.980 4.640 9.850 5.440 ;
        RECT  9.850 4.170 9.860 5.440 ;
        RECT  9.860 3.970 10.260 5.440 ;
        RECT  10.260 4.170 10.270 5.440 ;
        RECT  10.270 4.640 11.830 5.440 ;
        RECT  11.830 3.860 11.840 5.440 ;
        RECT  11.840 3.660 12.240 5.440 ;
        RECT  12.240 3.860 12.250 5.440 ;
        RECT  12.250 4.640 13.340 5.440 ;
        RECT  13.340 4.480 13.740 5.440 ;
        RECT  13.740 4.640 14.520 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.060 0.400 ;
        RECT  1.060 -0.400 1.460 0.560 ;
        RECT  1.460 -0.400 3.550 0.400 ;
        RECT  3.550 -0.400 3.560 0.730 ;
        RECT  3.560 -0.400 3.960 0.850 ;
        RECT  3.960 -0.400 3.970 0.730 ;
        RECT  3.970 -0.400 5.570 0.400 ;
        RECT  5.570 -0.400 5.830 1.530 ;
        RECT  5.830 1.290 7.350 1.530 ;
        RECT  7.350 1.290 7.590 1.840 ;
        RECT  7.590 1.440 7.750 1.840 ;
        RECT  5.830 -0.400 10.040 0.400 ;
        RECT  10.040 -0.400 10.440 1.280 ;
        RECT  10.440 -0.400 11.780 0.400 ;
        RECT  11.780 -0.400 11.790 0.690 ;
        RECT  11.790 -0.400 12.190 0.890 ;
        RECT  12.190 -0.400 12.200 0.690 ;
        RECT  12.200 -0.400 13.350 0.400 ;
        RECT  13.350 -0.400 13.750 0.560 ;
        RECT  13.750 -0.400 14.520 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.910 1.450 13.150 3.180 ;
        RECT  12.610 1.450 12.910 1.690 ;
        RECT  12.610 2.780 12.910 3.180 ;
        RECT  11.680 1.970 12.440 2.370 ;
        RECT  11.440 1.590 11.680 3.270 ;
        RECT  11.350 1.590 11.440 1.830 ;
        RECT  11.020 3.030 11.440 3.270 ;
        RECT  10.950 0.880 11.350 1.830 ;
        RECT  10.760 2.150 11.160 2.550 ;
        RECT  10.620 3.030 11.020 3.640 ;
        RECT  10.160 1.590 10.950 1.830 ;
        RECT  9.480 2.270 10.760 2.510 ;
        RECT  9.760 1.590 10.160 1.990 ;
        RECT  9.480 3.730 9.520 4.130 ;
        RECT  9.470 2.270 9.480 4.130 ;
        RECT  9.230 1.180 9.470 4.130 ;
        RECT  9.100 1.180 9.230 1.420 ;
        RECT  9.120 3.730 9.230 4.130 ;
        RECT  8.700 1.020 9.100 1.420 ;
        RECT  8.840 2.490 8.920 2.890 ;
        RECT  8.600 2.490 8.840 3.830 ;
        RECT  8.320 1.850 8.800 2.090 ;
        RECT  7.120 3.590 8.600 3.830 ;
        RECT  8.080 0.670 8.320 3.310 ;
        RECT  6.110 0.670 8.080 0.910 ;
        RECT  7.400 3.070 8.080 3.310 ;
        RECT  6.470 2.160 7.840 2.560 ;
        RECT  6.880 2.880 7.120 3.830 ;
        RECT  6.410 3.590 6.880 3.830 ;
        RECT  6.230 1.820 6.470 3.140 ;
        RECT  6.170 3.590 6.410 4.290 ;
        RECT  5.250 1.820 6.230 2.060 ;
        RECT  5.780 2.900 6.230 3.140 ;
        RECT  4.360 4.050 6.170 4.290 ;
        RECT  5.100 2.340 5.950 2.580 ;
        RECT  5.540 2.900 5.780 3.770 ;
        RECT  5.380 3.530 5.540 3.770 ;
        RECT  5.160 1.650 5.250 2.060 ;
        RECT  5.010 1.120 5.160 2.060 ;
        RECT  4.860 2.340 5.100 3.770 ;
        RECT  4.920 1.120 5.010 1.890 ;
        RECT  3.680 1.650 4.920 1.890 ;
        RECT  4.770 2.340 4.860 2.580 ;
        RECT  4.640 3.530 4.860 3.770 ;
        RECT  4.370 2.170 4.770 2.580 ;
        RECT  4.480 0.770 4.640 1.010 ;
        RECT  4.240 0.770 4.480 1.370 ;
        RECT  4.120 3.940 4.360 4.290 ;
        RECT  3.050 1.130 4.240 1.370 ;
        RECT  3.150 3.940 4.120 4.180 ;
        RECT  3.440 1.650 3.680 2.850 ;
        RECT  2.750 3.940 3.150 4.300 ;
        RECT  2.910 1.130 3.050 2.600 ;
        RECT  2.810 1.130 2.910 3.650 ;
        RECT  2.610 1.130 2.810 1.370 ;
        RECT  2.670 2.360 2.810 3.650 ;
        RECT  2.390 3.940 2.750 4.180 ;
        RECT  2.210 0.930 2.610 1.370 ;
        RECT  2.150 1.680 2.390 4.180 ;
        RECT  2.200 1.010 2.210 1.370 ;
        RECT  1.910 1.680 2.150 2.080 ;
        RECT  0.570 3.940 2.150 4.180 ;
        RECT  0.580 1.680 1.910 1.920 ;
        RECT  0.340 1.110 0.580 1.920 ;
        RECT  0.330 3.270 0.570 4.180 ;
        RECT  0.180 1.110 0.340 1.510 ;
        RECT  0.170 3.270 0.330 3.670 ;
    END
END DFFRX1

MACRO DFFNSRXL
    CLASS CORE ;
    FOREIGN DFFNSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.460 3.940 4.860 4.370 ;
        RECT  4.860 3.940 5.970 4.180 ;
        RECT  5.970 3.940 6.210 4.360 ;
        RECT  6.210 4.120 8.420 4.360 ;
        RECT  8.420 4.120 8.790 4.370 ;
        RECT  8.790 4.130 12.010 4.370 ;
        RECT  12.010 4.030 12.410 4.370 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.040 1.770 6.560 2.190 ;
        RECT  6.560 1.780 6.780 2.180 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.720 1.830 14.880 2.090 ;
        RECT  14.880 1.390 15.120 3.210 ;
        RECT  15.120 1.390 15.280 1.790 ;
        RECT  15.120 2.810 15.340 3.210 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.590 1.390 16.610 1.790 ;
        RECT  16.590 2.900 16.700 3.300 ;
        RECT  16.700 2.390 16.710 3.300 ;
        RECT  16.610 1.390 16.710 1.820 ;
        RECT  16.710 1.390 16.950 3.300 ;
        RECT  16.950 2.390 16.960 3.300 ;
        RECT  16.960 2.900 16.990 3.300 ;
        RECT  16.950 1.390 16.990 1.950 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.390 1.610 2.650 ;
        RECT  1.610 2.100 1.780 2.650 ;
        RECT  1.780 2.100 2.010 2.640 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.720 1.740 1.210 2.140 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 4.480 1.390 5.440 ;
        RECT  1.390 4.640 3.680 5.440 ;
        RECT  3.680 4.480 4.080 5.440 ;
        RECT  4.080 4.640 5.290 5.440 ;
        RECT  5.290 4.480 5.690 5.440 ;
        RECT  9.100 3.510 9.500 3.850 ;
        RECT  9.500 3.610 11.310 3.850 ;
        RECT  11.310 3.460 11.550 3.850 ;
        RECT  5.690 4.640 12.710 5.440 ;
        RECT  11.550 3.460 12.710 3.700 ;
        RECT  12.710 3.460 12.950 5.440 ;
        RECT  12.950 4.640 13.890 5.440 ;
        RECT  13.890 3.650 13.900 5.440 ;
        RECT  13.900 3.450 14.300 5.440 ;
        RECT  14.300 3.650 14.310 5.440 ;
        RECT  14.310 4.640 15.750 5.440 ;
        RECT  15.750 4.480 16.150 5.440 ;
        RECT  16.150 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.250 0.400 ;
        RECT  1.250 -0.400 1.650 0.560 ;
        RECT  1.650 -0.400 3.890 0.400 ;
        RECT  3.890 -0.400 3.900 0.730 ;
        RECT  3.900 -0.400 4.300 0.930 ;
        RECT  4.300 -0.400 4.310 0.730 ;
        RECT  4.310 -0.400 6.940 0.400 ;
        RECT  6.940 -0.400 6.950 0.730 ;
        RECT  6.950 -0.400 7.350 0.850 ;
        RECT  7.350 -0.400 7.360 0.730 ;
        RECT  7.360 -0.400 9.190 0.400 ;
        RECT  9.190 -0.400 9.200 0.750 ;
        RECT  9.200 -0.400 9.600 0.870 ;
        RECT  9.600 -0.400 9.610 0.750 ;
        RECT  9.610 -0.400 11.770 0.400 ;
        RECT  11.770 -0.400 12.170 0.560 ;
        RECT  12.170 -0.400 15.770 0.400 ;
        RECT  15.770 -0.400 16.170 0.560 ;
        RECT  16.170 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.180 2.220 16.340 2.620 ;
        RECT  15.940 0.860 16.180 3.980 ;
        RECT  15.280 0.860 15.940 1.100 ;
        RECT  15.280 3.740 15.940 3.980 ;
        RECT  15.040 0.740 15.280 1.100 ;
        RECT  14.880 3.740 15.280 4.140 ;
        RECT  14.880 0.740 15.040 0.980 ;
        RECT  14.140 2.460 14.600 2.860 ;
        RECT  13.900 1.480 14.140 3.170 ;
        RECT  13.300 1.480 13.900 1.720 ;
        RECT  11.840 2.930 13.900 3.170 ;
        RECT  12.860 1.990 13.260 2.390 ;
        RECT  11.060 1.990 12.860 2.230 ;
        RECT  11.440 2.770 11.840 3.170 ;
        RECT  10.280 0.730 11.340 0.970 ;
        RECT  11.020 1.290 11.060 2.230 ;
        RECT  10.780 1.290 11.020 3.330 ;
        RECT  10.640 1.290 10.780 1.530 ;
        RECT  10.400 3.090 10.780 3.330 ;
        RECT  10.280 2.520 10.500 2.760 ;
        RECT  10.040 0.730 10.280 2.760 ;
        RECT  8.660 1.150 10.040 1.390 ;
        RECT  9.930 2.520 10.040 2.760 ;
        RECT  9.690 2.520 9.930 3.130 ;
        RECT  7.980 1.850 9.740 2.090 ;
        RECT  8.660 2.890 9.690 3.130 ;
        RECT  8.030 2.370 9.020 2.610 ;
        RECT  8.500 1.150 8.660 1.570 ;
        RECT  8.420 2.890 8.660 3.830 ;
        RECT  8.260 0.670 8.500 1.570 ;
        RECT  7.790 2.370 8.030 3.840 ;
        RECT  7.740 1.130 7.980 2.090 ;
        RECT  6.730 3.600 7.790 3.840 ;
        RECT  5.840 1.130 7.740 1.370 ;
        RECT  7.460 2.430 7.500 3.320 ;
        RECT  7.220 1.650 7.460 3.320 ;
        RECT  7.050 1.650 7.220 1.890 ;
        RECT  7.010 2.900 7.220 3.320 ;
        RECT  6.280 2.900 7.010 3.140 ;
        RECT  6.490 3.420 6.730 3.840 ;
        RECT  3.100 3.420 6.490 3.660 ;
        RECT  6.040 2.510 6.280 3.140 ;
        RECT  5.760 1.100 5.840 1.500 ;
        RECT  5.520 1.100 5.760 3.140 ;
        RECT  5.440 1.100 5.520 1.500 ;
        RECT  3.780 2.900 5.520 3.140 ;
        RECT  5.150 1.790 5.240 2.200 ;
        RECT  4.910 1.230 5.150 2.200 ;
        RECT  2.990 1.230 4.910 1.470 ;
        RECT  3.380 2.740 3.780 3.140 ;
        RECT  3.100 1.750 3.230 2.150 ;
        RECT  2.860 1.750 3.100 4.180 ;
        RECT  2.590 1.070 2.990 1.470 ;
        RECT  2.420 3.940 2.860 4.180 ;
        RECT  2.580 1.230 2.590 1.470 ;
        RECT  2.340 1.230 2.580 3.630 ;
        RECT  2.020 3.940 2.420 4.360 ;
        RECT  0.500 3.940 2.020 4.180 ;
        RECT  0.480 1.260 0.760 1.500 ;
        RECT  0.480 3.040 0.500 4.180 ;
        RECT  0.260 1.260 0.480 4.180 ;
        RECT  0.240 1.260 0.260 3.360 ;
    END
END DFFNSRXL

MACRO DFFNSRX4
    CLASS CORE ;
    FOREIGN DFFNSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNSRXL ;
    SIZE 23.100 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.100 3.990 4.500 4.360 ;
        RECT  4.500 4.120 8.040 4.360 ;
        RECT  8.040 3.940 8.460 4.360 ;
        RECT  8.460 3.940 12.990 4.180 ;
        RECT  12.990 3.940 13.380 4.350 ;
        RECT  13.380 3.940 13.690 4.340 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.050 2.380 6.520 2.810 ;
        RECT  6.520 2.400 6.590 2.800 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  19.910 1.820 20.080 3.220 ;
        RECT  20.080 1.590 20.090 3.220 ;
        RECT  20.090 1.390 20.350 3.220 ;
        RECT  20.350 1.390 20.490 3.150 ;
        RECT  20.490 1.590 20.500 2.950 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.230 1.820 21.400 3.220 ;
        RECT  21.400 1.590 21.410 3.220 ;
        RECT  21.410 1.390 21.670 3.220 ;
        RECT  21.670 1.390 21.810 3.160 ;
        RECT  21.810 1.590 21.820 3.150 ;
        RECT  21.820 2.750 22.010 3.150 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.240 2.530 1.400 2.930 ;
        RECT  1.400 2.530 1.520 3.190 ;
        RECT  1.520 2.530 1.640 3.210 ;
        RECT  1.640 2.950 1.780 3.210 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 1.820 0.690 2.210 ;
        RECT  0.690 1.800 1.090 2.210 ;
        RECT  1.090 1.820 1.140 2.210 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.980 5.440 ;
        RECT  0.980 4.480 1.380 5.440 ;
        RECT  1.380 4.640 3.430 5.440 ;
        RECT  3.430 4.480 3.830 5.440 ;
        RECT  3.830 4.640 8.950 5.440 ;
        RECT  8.950 4.480 9.350 5.440 ;
        RECT  9.350 4.640 11.510 5.440 ;
        RECT  11.510 4.480 11.910 5.440 ;
        RECT  11.910 4.640 14.630 5.440 ;
        RECT  14.630 3.110 15.030 5.440 ;
        RECT  15.030 4.640 16.600 5.440 ;
        RECT  16.600 3.810 16.610 5.440 ;
        RECT  16.610 3.610 17.010 5.440 ;
        RECT  17.010 3.810 17.020 5.440 ;
        RECT  17.020 4.640 19.420 5.440 ;
        RECT  19.420 4.210 19.430 5.440 ;
        RECT  19.430 4.010 19.830 5.440 ;
        RECT  19.830 4.210 19.840 5.440 ;
        RECT  19.840 4.640 20.860 5.440 ;
        RECT  20.860 4.210 20.870 5.440 ;
        RECT  20.870 4.010 21.270 5.440 ;
        RECT  21.270 4.210 21.280 5.440 ;
        RECT  21.280 4.640 22.270 5.440 ;
        RECT  22.270 4.210 22.280 5.440 ;
        RECT  22.280 4.010 22.680 5.440 ;
        RECT  22.680 4.210 22.690 5.440 ;
        RECT  22.690 4.640 23.100 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.040 0.400 ;
        RECT  1.040 -0.400 1.440 0.560 ;
        RECT  1.440 -0.400 3.300 0.400 ;
        RECT  3.300 -0.400 3.310 0.730 ;
        RECT  3.310 -0.400 3.710 0.850 ;
        RECT  3.710 -0.400 3.720 0.730 ;
        RECT  3.720 -0.400 6.720 0.400 ;
        RECT  6.720 -0.400 6.730 0.800 ;
        RECT  6.730 -0.400 7.130 0.920 ;
        RECT  7.130 -0.400 7.140 0.800 ;
        RECT  7.140 -0.400 8.780 0.400 ;
        RECT  8.780 -0.400 8.790 0.860 ;
        RECT  8.790 -0.400 9.190 0.980 ;
        RECT  9.190 -0.400 9.200 0.860 ;
        RECT  9.200 -0.400 11.340 0.400 ;
        RECT  11.340 -0.400 11.350 0.820 ;
        RECT  11.350 -0.400 11.750 0.940 ;
        RECT  11.750 -0.400 11.760 0.820 ;
        RECT  11.760 -0.400 14.280 0.400 ;
        RECT  14.280 -0.400 14.290 1.100 ;
        RECT  14.290 -0.400 14.690 1.220 ;
        RECT  14.690 -0.400 14.700 1.100 ;
        RECT  14.700 -0.400 19.470 0.400 ;
        RECT  19.470 -0.400 19.480 0.910 ;
        RECT  19.480 -0.400 19.880 1.110 ;
        RECT  19.880 -0.400 19.890 0.910 ;
        RECT  19.890 -0.400 20.750 0.400 ;
        RECT  20.750 -0.400 20.760 0.910 ;
        RECT  20.760 -0.400 21.160 1.110 ;
        RECT  21.160 -0.400 21.170 0.910 ;
        RECT  21.170 -0.400 22.070 0.400 ;
        RECT  22.070 -0.400 22.080 0.910 ;
        RECT  22.080 -0.400 22.480 1.110 ;
        RECT  22.480 -0.400 22.490 0.910 ;
        RECT  22.490 -0.400 23.100 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  22.290 2.180 22.530 3.730 ;
        RECT  19.640 3.490 22.290 3.730 ;
        RECT  19.400 1.550 19.640 3.730 ;
        RECT  18.980 1.550 19.400 1.790 ;
        RECT  18.610 3.330 19.400 3.730 ;
        RECT  18.720 2.130 19.120 2.530 ;
        RECT  18.740 1.390 18.980 1.790 ;
        RECT  18.410 2.140 18.720 2.530 ;
        RECT  18.410 0.720 18.490 0.960 ;
        RECT  18.090 0.680 18.410 0.960 ;
        RECT  18.230 1.370 18.410 3.020 ;
        RECT  18.170 1.370 18.230 3.640 ;
        RECT  17.730 1.370 18.170 1.610 ;
        RECT  17.990 2.780 18.170 3.640 ;
        RECT  16.970 0.680 18.090 0.920 ;
        RECT  17.830 3.080 17.990 3.640 ;
        RECT  17.650 1.890 17.890 2.290 ;
        RECT  15.790 3.080 17.830 3.320 ;
        RECT  17.330 1.200 17.730 1.610 ;
        RECT  15.990 1.990 17.650 2.230 ;
        RECT  16.210 1.370 17.330 1.610 ;
        RECT  16.570 0.680 16.970 1.080 ;
        RECT  15.450 0.680 16.570 0.920 ;
        RECT  15.810 1.240 16.210 1.610 ;
        RECT  15.590 1.910 15.990 2.310 ;
        RECT  15.630 3.080 15.790 3.630 ;
        RECT  15.390 2.590 15.630 3.630 ;
        RECT  13.300 2.070 15.590 2.310 ;
        RECT  15.290 0.680 15.450 1.500 ;
        RECT  14.270 2.590 15.390 2.830 ;
        RECT  15.210 0.680 15.290 1.740 ;
        RECT  15.050 1.100 15.210 1.740 ;
        RECT  13.850 1.500 15.050 1.740 ;
        RECT  14.110 3.420 14.350 4.370 ;
        RECT  14.030 2.590 14.270 3.140 ;
        RECT  7.860 3.420 14.110 3.660 ;
        RECT  13.870 2.870 14.030 3.140 ;
        RECT  12.180 2.900 13.870 3.140 ;
        RECT  13.610 0.790 13.850 1.740 ;
        RECT  13.060 0.830 13.300 2.310 ;
        RECT  12.690 0.830 13.060 1.070 ;
        RECT  12.870 1.920 13.060 2.310 ;
        RECT  12.470 1.920 12.870 2.620 ;
        RECT  12.340 1.400 12.770 1.640 ;
        RECT  10.910 1.920 12.470 2.160 ;
        RECT  12.100 1.230 12.340 1.640 ;
        RECT  11.940 2.440 12.180 3.140 ;
        RECT  11.070 1.230 12.100 1.470 ;
        RECT  11.780 2.440 11.940 2.680 ;
        RECT  10.830 0.670 11.070 1.470 ;
        RECT  10.670 1.750 10.910 3.140 ;
        RECT  9.750 0.670 10.830 0.910 ;
        RECT  10.390 1.750 10.670 1.990 ;
        RECT  10.230 2.900 10.670 3.140 ;
        RECT  10.150 1.190 10.390 1.990 ;
        RECT  9.750 2.270 10.390 2.510 ;
        RECT  9.510 0.670 9.750 2.910 ;
        RECT  8.210 1.260 9.510 1.500 ;
        RECT  8.540 2.670 9.510 2.910 ;
        RECT  8.990 1.780 9.230 2.180 ;
        RECT  7.690 1.860 8.990 2.100 ;
        RECT  8.140 2.670 8.540 3.140 ;
        RECT  7.970 0.680 8.210 1.580 ;
        RECT  7.540 0.680 7.970 0.920 ;
        RECT  7.620 3.080 7.860 3.660 ;
        RECT  7.450 1.200 7.690 2.100 ;
        RECT  7.170 3.080 7.620 3.320 ;
        RECT  6.490 1.200 7.450 1.440 ;
        RECT  5.040 3.600 7.340 3.840 ;
        RECT  6.930 1.720 7.170 3.320 ;
        RECT  6.770 1.720 6.930 1.960 ;
        RECT  5.730 3.080 6.930 3.320 ;
        RECT  6.250 1.200 6.490 1.990 ;
        RECT  5.290 1.750 6.250 1.990 ;
        RECT  5.730 0.670 5.970 1.470 ;
        RECT  4.450 0.670 5.730 0.910 ;
        RECT  5.490 2.370 5.730 3.320 ;
        RECT  5.210 1.190 5.290 1.990 ;
        RECT  4.970 1.190 5.210 3.100 ;
        RECT  4.800 3.470 5.040 3.840 ;
        RECT  4.890 1.190 4.970 1.430 ;
        RECT  4.750 2.860 4.970 3.100 ;
        RECT  3.010 3.470 4.800 3.710 ;
        RECT  4.350 2.860 4.750 3.190 ;
        RECT  4.450 1.710 4.690 2.140 ;
        RECT  4.210 0.670 4.450 1.370 ;
        RECT  3.910 1.710 4.450 1.950 ;
        RECT  3.530 2.860 4.350 3.100 ;
        RECT  3.670 1.220 3.910 1.950 ;
        RECT  2.290 1.220 3.670 1.460 ;
        RECT  3.290 2.300 3.530 3.100 ;
        RECT  2.770 1.740 3.010 4.170 ;
        RECT  2.570 1.740 2.770 2.140 ;
        RECT  2.340 3.930 2.770 4.170 ;
        RECT  2.290 2.420 2.490 3.520 ;
        RECT  1.940 3.930 2.340 4.370 ;
        RECT  2.250 1.220 2.290 3.520 ;
        RECT  2.050 1.220 2.250 2.660 ;
        RECT  0.570 3.930 1.940 4.170 ;
        RECT  0.400 1.090 0.570 1.490 ;
        RECT  0.400 3.120 0.570 4.170 ;
        RECT  0.170 1.090 0.400 4.170 ;
        RECT  0.160 1.250 0.170 4.170 ;
    END
END DFFNSRX4

MACRO DFFNSRX2
    CLASS CORE ;
    FOREIGN DFFNSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNSRXL ;
    SIZE 17.820 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.540 3.940 4.940 4.370 ;
        RECT  4.940 3.940 5.970 4.180 ;
        RECT  5.970 3.940 6.210 4.360 ;
        RECT  6.210 4.120 8.420 4.360 ;
        RECT  8.420 4.120 8.790 4.370 ;
        RECT  8.790 4.130 12.010 4.370 ;
        RECT  12.010 4.030 12.410 4.370 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.140 1.770 6.790 2.190 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.380 2.950 15.500 3.210 ;
        RECT  15.500 2.640 15.540 3.210 ;
        RECT  15.540 1.160 15.740 3.210 ;
        RECT  15.740 1.160 15.780 3.050 ;
        RECT  15.780 1.160 16.130 1.560 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.700 2.950 16.810 3.210 ;
        RECT  16.810 2.950 17.150 3.220 ;
        RECT  17.150 2.950 17.410 4.160 ;
        RECT  17.250 0.950 17.410 1.350 ;
        RECT  17.410 0.950 17.550 4.160 ;
        RECT  17.550 0.950 17.650 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 2.940 1.870 3.360 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.770 2.230 1.210 2.660 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.110 5.440 ;
        RECT  1.110 4.480 1.510 5.440 ;
        RECT  1.510 4.640 3.860 5.440 ;
        RECT  3.860 4.480 4.260 5.440 ;
        RECT  4.260 4.640 5.290 5.440 ;
        RECT  5.290 4.480 5.690 5.440 ;
        RECT  9.100 3.510 9.500 3.850 ;
        RECT  9.500 3.610 11.310 3.850 ;
        RECT  11.310 3.460 11.550 3.850 ;
        RECT  5.690 4.640 12.710 5.440 ;
        RECT  11.550 3.460 12.710 3.700 ;
        RECT  12.710 3.460 12.950 5.440 ;
        RECT  12.950 4.640 13.830 5.440 ;
        RECT  13.830 3.730 13.840 5.440 ;
        RECT  13.840 3.530 14.240 5.440 ;
        RECT  14.240 3.730 14.250 5.440 ;
        RECT  14.250 4.640 16.330 5.440 ;
        RECT  16.330 4.150 16.730 5.440 ;
        RECT  16.730 4.640 17.820 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.120 0.400 ;
        RECT  1.120 -0.400 1.130 1.300 ;
        RECT  1.130 -0.400 1.530 1.420 ;
        RECT  1.530 -0.400 1.540 1.300 ;
        RECT  1.540 -0.400 3.890 0.400 ;
        RECT  3.890 -0.400 3.900 0.730 ;
        RECT  3.900 -0.400 4.300 0.850 ;
        RECT  4.300 -0.400 4.310 0.730 ;
        RECT  4.310 -0.400 6.950 0.400 ;
        RECT  6.950 -0.400 7.350 0.850 ;
        RECT  7.350 -0.400 9.190 0.400 ;
        RECT  9.190 -0.400 9.200 0.750 ;
        RECT  9.200 -0.400 9.600 0.870 ;
        RECT  9.600 -0.400 9.610 0.750 ;
        RECT  9.610 -0.400 11.770 0.400 ;
        RECT  11.770 -0.400 12.170 0.560 ;
        RECT  12.170 -0.400 14.930 0.400 ;
        RECT  14.930 -0.400 15.330 0.560 ;
        RECT  15.330 -0.400 16.480 0.400 ;
        RECT  16.480 -0.400 16.490 1.220 ;
        RECT  16.490 -0.400 16.890 1.710 ;
        RECT  16.890 -0.400 16.900 1.220 ;
        RECT  16.900 -0.400 17.820 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.710 2.240 17.110 2.640 ;
        RECT  16.340 2.400 16.710 2.640 ;
        RECT  16.100 2.400 16.340 3.730 ;
        RECT  15.070 3.490 16.100 3.730 ;
        RECT  15.020 1.300 15.260 1.700 ;
        RECT  15.020 3.490 15.070 3.890 ;
        RECT  14.780 1.300 15.020 3.890 ;
        RECT  14.670 3.490 14.780 3.890 ;
        RECT  14.420 0.750 14.500 1.150 ;
        RECT  13.740 2.270 14.500 2.670 ;
        RECT  14.100 0.740 14.420 1.150 ;
        RECT  12.980 0.740 14.100 0.980 ;
        RECT  13.500 1.270 13.740 3.170 ;
        RECT  13.340 1.270 13.500 1.510 ;
        RECT  11.810 2.930 13.500 3.170 ;
        RECT  12.820 1.790 13.220 2.190 ;
        RECT  12.660 0.740 12.980 1.150 ;
        RECT  11.060 1.850 12.820 2.090 ;
        RECT  12.580 0.750 12.660 1.150 ;
        RECT  11.570 2.610 11.810 3.170 ;
        RECT  11.400 2.610 11.570 2.850 ;
        RECT  10.280 0.730 11.340 0.970 ;
        RECT  11.020 1.330 11.060 2.090 ;
        RECT  10.780 1.330 11.020 3.330 ;
        RECT  10.640 1.330 10.780 1.570 ;
        RECT  10.400 3.090 10.780 3.330 ;
        RECT  10.280 2.520 10.500 2.760 ;
        RECT  10.040 0.730 10.280 2.760 ;
        RECT  8.660 1.150 10.040 1.390 ;
        RECT  9.930 2.520 10.040 2.760 ;
        RECT  9.690 2.520 9.930 3.130 ;
        RECT  9.340 1.850 9.740 2.140 ;
        RECT  8.660 2.890 9.690 3.130 ;
        RECT  7.980 1.850 9.340 2.090 ;
        RECT  8.030 2.370 9.020 2.610 ;
        RECT  8.500 1.150 8.660 1.570 ;
        RECT  8.420 2.890 8.660 3.830 ;
        RECT  8.260 0.670 8.500 1.570 ;
        RECT  7.790 2.370 8.030 3.840 ;
        RECT  7.740 1.130 7.980 2.090 ;
        RECT  6.730 3.600 7.790 3.840 ;
        RECT  6.570 1.130 7.740 1.370 ;
        RECT  7.460 2.430 7.500 3.140 ;
        RECT  7.410 1.650 7.460 3.140 ;
        RECT  7.220 1.650 7.410 3.360 ;
        RECT  7.060 1.650 7.220 1.890 ;
        RECT  7.010 2.900 7.220 3.360 ;
        RECT  6.280 2.900 7.010 3.140 ;
        RECT  6.490 3.420 6.730 3.840 ;
        RECT  6.330 1.130 6.570 1.430 ;
        RECT  3.560 3.420 6.490 3.660 ;
        RECT  5.760 1.190 6.330 1.430 ;
        RECT  6.040 2.510 6.280 3.140 ;
        RECT  5.520 1.190 5.760 3.140 ;
        RECT  5.440 1.190 5.520 1.430 ;
        RECT  4.080 2.900 5.520 3.140 ;
        RECT  5.000 1.740 5.240 2.190 ;
        RECT  4.100 1.740 5.000 1.980 ;
        RECT  3.860 1.210 4.100 1.980 ;
        RECT  3.840 2.490 4.080 3.140 ;
        RECT  2.920 1.210 3.860 1.450 ;
        RECT  3.320 1.740 3.560 4.370 ;
        RECT  3.180 1.740 3.320 2.140 ;
        RECT  2.470 4.130 3.320 4.370 ;
        RECT  3.000 3.450 3.040 3.850 ;
        RECT  2.900 2.430 3.000 3.850 ;
        RECT  2.900 1.130 2.920 1.450 ;
        RECT  2.760 1.130 2.900 3.850 ;
        RECT  2.660 1.130 2.760 2.670 ;
        RECT  2.520 1.130 2.660 1.370 ;
        RECT  2.380 2.950 2.470 4.370 ;
        RECT  2.230 1.700 2.380 4.370 ;
        RECT  2.140 1.700 2.230 3.270 ;
        RECT  0.650 1.700 2.140 1.940 ;
        RECT  0.500 3.400 0.680 3.800 ;
        RECT  0.500 1.330 0.650 1.940 ;
        RECT  0.260 1.330 0.500 3.800 ;
        RECT  0.250 1.330 0.260 1.730 ;
    END
END DFFNSRX2

MACRO DFFNSRX1
    CLASS CORE ;
    FOREIGN DFFNSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNSRXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.540 4.130 4.670 4.370 ;
        RECT  4.670 3.940 4.940 4.370 ;
        RECT  4.940 3.940 5.970 4.180 ;
        RECT  5.970 3.940 6.210 4.360 ;
        RECT  6.210 4.120 8.420 4.360 ;
        RECT  8.420 4.120 8.790 4.370 ;
        RECT  8.790 4.130 12.010 4.370 ;
        RECT  12.010 4.030 12.410 4.370 ;
        END
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.140 1.770 6.690 2.190 ;
        RECT  6.690 1.780 6.780 2.180 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.180 0.740 14.420 3.090 ;
        RECT  14.420 0.740 14.720 0.980 ;
        RECT  14.720 0.710 14.970 0.980 ;
        RECT  14.970 0.710 14.980 0.970 ;
        RECT  14.420 2.850 15.100 3.090 ;
        RECT  14.980 0.730 15.160 0.970 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.590 2.970 16.710 3.370 ;
        RECT  16.700 2.390 16.710 2.650 ;
        RECT  16.590 1.320 16.710 1.960 ;
        RECT  16.710 1.320 16.950 3.370 ;
        RECT  16.950 2.390 16.960 2.650 ;
        RECT  16.950 2.970 16.990 3.370 ;
        RECT  16.950 1.320 16.990 1.960 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.500 1.950 1.520 2.350 ;
        RECT  1.520 1.830 1.780 2.350 ;
        RECT  1.780 1.950 1.900 2.350 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.800 2.650 0.860 3.070 ;
        RECT  0.860 2.390 1.120 3.070 ;
        RECT  1.120 2.650 1.200 3.070 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.110 5.440 ;
        RECT  1.110 4.480 1.510 5.440 ;
        RECT  1.510 4.640 3.860 5.440 ;
        RECT  3.860 4.480 4.260 5.440 ;
        RECT  4.260 4.640 5.290 5.440 ;
        RECT  5.290 4.480 5.690 5.440 ;
        RECT  9.100 3.510 9.260 3.750 ;
        RECT  9.260 3.510 9.500 3.850 ;
        RECT  9.500 3.610 11.310 3.850 ;
        RECT  11.310 3.460 11.550 3.850 ;
        RECT  5.690 4.640 12.710 5.440 ;
        RECT  11.550 3.460 12.710 3.700 ;
        RECT  12.710 3.460 12.950 5.440 ;
        RECT  12.950 4.640 13.890 5.440 ;
        RECT  13.890 4.050 13.900 5.440 ;
        RECT  13.900 3.930 14.300 5.440 ;
        RECT  14.300 4.050 14.310 5.440 ;
        RECT  14.310 4.640 15.520 5.440 ;
        RECT  15.520 4.480 15.920 5.440 ;
        RECT  15.920 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.170 0.400 ;
        RECT  1.170 -0.400 1.180 1.400 ;
        RECT  1.180 -0.400 1.580 1.520 ;
        RECT  1.580 -0.400 1.590 1.400 ;
        RECT  1.590 -0.400 3.890 0.400 ;
        RECT  3.890 -0.400 3.900 0.730 ;
        RECT  3.900 -0.400 4.300 0.850 ;
        RECT  4.300 -0.400 4.310 0.730 ;
        RECT  4.310 -0.400 6.940 0.400 ;
        RECT  6.940 -0.400 6.950 0.730 ;
        RECT  6.950 -0.400 7.350 0.850 ;
        RECT  7.350 -0.400 7.360 0.730 ;
        RECT  7.360 -0.400 9.190 0.400 ;
        RECT  9.190 -0.400 9.200 0.930 ;
        RECT  9.200 -0.400 9.600 1.050 ;
        RECT  9.600 -0.400 9.610 0.930 ;
        RECT  9.610 -0.400 11.760 0.400 ;
        RECT  11.760 -0.400 12.160 0.560 ;
        RECT  12.160 -0.400 15.650 0.400 ;
        RECT  15.650 -0.400 15.660 1.070 ;
        RECT  15.660 -0.400 16.060 1.270 ;
        RECT  16.060 -0.400 16.070 1.070 ;
        RECT  16.070 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.180 2.180 16.340 2.580 ;
        RECT  15.940 1.550 16.180 4.170 ;
        RECT  15.100 1.550 15.940 1.790 ;
        RECT  15.040 3.930 15.940 4.170 ;
        RECT  15.420 2.170 15.660 3.610 ;
        RECT  15.300 2.170 15.420 2.570 ;
        RECT  13.800 3.370 15.420 3.610 ;
        RECT  14.700 1.390 15.100 1.790 ;
        RECT  14.640 3.930 15.040 4.330 ;
        RECT  13.560 1.490 13.800 3.610 ;
        RECT  13.540 1.490 13.560 1.730 ;
        RECT  11.840 2.930 13.560 3.170 ;
        RECT  13.140 1.330 13.540 1.730 ;
        RECT  12.860 2.160 13.260 2.560 ;
        RECT  11.060 2.160 12.860 2.400 ;
        RECT  11.600 2.680 11.840 3.170 ;
        RECT  11.430 2.680 11.600 2.920 ;
        RECT  10.260 0.730 11.240 0.970 ;
        RECT  11.020 1.300 11.060 2.400 ;
        RECT  10.780 1.300 11.020 3.330 ;
        RECT  10.540 1.300 10.780 1.540 ;
        RECT  10.400 3.090 10.780 3.330 ;
        RECT  10.260 2.520 10.500 2.760 ;
        RECT  10.020 0.730 10.260 2.760 ;
        RECT  9.920 0.730 10.020 1.570 ;
        RECT  9.930 2.520 10.020 2.760 ;
        RECT  9.690 2.520 9.930 3.130 ;
        RECT  8.500 1.330 9.920 1.570 ;
        RECT  9.340 1.850 9.740 2.110 ;
        RECT  8.660 2.890 9.690 3.130 ;
        RECT  7.980 1.850 9.340 2.090 ;
        RECT  8.030 2.370 9.020 2.610 ;
        RECT  8.420 2.890 8.660 3.830 ;
        RECT  8.260 0.670 8.500 1.570 ;
        RECT  7.790 2.370 8.030 3.840 ;
        RECT  7.740 1.130 7.980 2.090 ;
        RECT  6.730 3.600 7.790 3.840 ;
        RECT  6.570 1.130 7.740 1.370 ;
        RECT  7.460 2.430 7.500 3.320 ;
        RECT  7.220 1.650 7.460 3.320 ;
        RECT  7.050 1.650 7.220 1.890 ;
        RECT  7.010 2.900 7.220 3.320 ;
        RECT  6.280 2.900 7.010 3.140 ;
        RECT  6.490 3.420 6.730 3.840 ;
        RECT  6.330 1.130 6.570 1.410 ;
        RECT  3.560 3.420 6.490 3.660 ;
        RECT  5.760 1.170 6.330 1.410 ;
        RECT  6.040 2.510 6.280 3.140 ;
        RECT  5.520 1.170 5.760 3.140 ;
        RECT  5.440 1.170 5.520 1.410 ;
        RECT  4.080 2.900 5.520 3.140 ;
        RECT  5.000 1.740 5.240 2.190 ;
        RECT  4.100 1.740 5.000 1.980 ;
        RECT  3.860 1.130 4.100 1.980 ;
        RECT  3.840 2.610 4.080 3.140 ;
        RECT  2.900 1.130 3.860 1.370 ;
        RECT  3.320 1.740 3.560 4.360 ;
        RECT  3.180 1.740 3.320 2.140 ;
        RECT  2.480 4.120 3.320 4.360 ;
        RECT  3.000 3.440 3.040 3.840 ;
        RECT  2.900 2.420 3.000 3.840 ;
        RECT  2.760 1.130 2.900 3.840 ;
        RECT  2.660 1.130 2.760 2.660 ;
        RECT  2.600 1.330 2.660 1.730 ;
        RECT  2.470 3.250 2.480 4.360 ;
        RECT  2.240 2.940 2.470 4.360 ;
        RECT  2.230 2.940 2.240 3.630 ;
        RECT  0.690 3.390 2.230 3.630 ;
        RECT  0.500 3.390 0.690 3.790 ;
        RECT  0.500 1.410 0.630 1.650 ;
        RECT  0.260 1.410 0.500 3.790 ;
        RECT  0.230 1.410 0.260 1.650 ;
    END
END DFFNSRX1

MACRO DFFNSXL
    CLASS CORE ;
    FOREIGN DFFNSXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  10.100 4.070 10.360 4.330 ;
        RECT  10.360 4.070 10.450 4.310 ;
        RECT  10.450 3.740 10.690 4.310 ;
        RECT  10.690 3.740 10.850 4.140 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.890 0.700 12.050 0.940 ;
        RECT  11.830 3.520 12.080 3.950 ;
        RECT  12.080 3.510 12.230 3.950 ;
        RECT  12.050 0.700 12.290 1.100 ;
        RECT  12.230 3.510 12.340 3.770 ;
        RECT  12.290 0.860 12.650 1.100 ;
        RECT  12.340 3.520 12.790 3.760 ;
        RECT  12.650 0.860 12.790 1.280 ;
        RECT  12.790 0.860 13.030 3.760 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.360 1.280 13.660 3.570 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.640 2.090 ;
        RECT  1.640 1.830 1.650 2.230 ;
        RECT  1.650 1.830 2.050 2.300 ;
        RECT  2.050 1.830 2.060 2.230 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.840 2.370 0.960 2.770 ;
        RECT  0.960 2.360 1.290 2.780 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.360 5.440 ;
        RECT  1.360 4.480 1.760 5.440 ;
        RECT  1.760 4.640 4.060 5.440 ;
        RECT  4.060 4.480 4.460 5.440 ;
        RECT  4.460 4.640 5.580 5.440 ;
        RECT  5.580 4.310 5.590 5.440 ;
        RECT  5.590 4.190 5.990 5.440 ;
        RECT  5.990 4.310 6.000 5.440 ;
        RECT  6.000 4.640 6.900 5.440 ;
        RECT  6.900 4.040 6.910 5.440 ;
        RECT  6.910 3.840 7.310 5.440 ;
        RECT  7.310 4.040 7.320 5.440 ;
        RECT  7.320 4.640 9.300 5.440 ;
        RECT  9.300 4.210 9.310 5.440 ;
        RECT  9.310 4.010 9.710 5.440 ;
        RECT  9.710 4.210 9.720 5.440 ;
        RECT  9.720 4.640 11.150 5.440 ;
        RECT  11.150 3.730 11.390 5.440 ;
        RECT  11.390 4.640 12.620 5.440 ;
        RECT  12.620 4.480 13.020 5.440 ;
        RECT  13.020 4.640 13.860 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.380 0.400 ;
        RECT  1.380 -0.400 1.390 1.420 ;
        RECT  1.390 -0.400 1.790 1.540 ;
        RECT  1.790 -0.400 1.800 1.420 ;
        RECT  1.800 -0.400 4.000 0.400 ;
        RECT  4.000 -0.400 4.010 0.750 ;
        RECT  4.010 -0.400 4.410 0.870 ;
        RECT  4.410 -0.400 4.420 0.750 ;
        RECT  4.420 -0.400 6.660 0.400 ;
        RECT  6.660 -0.400 6.670 0.750 ;
        RECT  6.670 -0.400 7.070 0.870 ;
        RECT  7.070 -0.400 7.080 0.750 ;
        RECT  7.080 -0.400 8.930 0.400 ;
        RECT  8.930 -0.400 9.330 0.560 ;
        RECT  9.330 -0.400 11.000 0.400 ;
        RECT  11.000 -0.400 11.010 0.850 ;
        RECT  11.010 -0.400 11.410 1.050 ;
        RECT  11.410 -0.400 11.420 0.850 ;
        RECT  11.420 -0.400 12.620 0.400 ;
        RECT  12.620 -0.400 13.020 0.560 ;
        RECT  13.020 -0.400 13.860 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.300 1.960 12.510 2.370 ;
        RECT  12.290 1.500 12.300 2.370 ;
        RECT  12.050 1.380 12.290 3.210 ;
        RECT  12.040 1.380 12.050 2.110 ;
        RECT  11.890 2.810 12.050 3.210 ;
        RECT  11.890 1.380 12.040 1.780 ;
        RECT  11.450 2.020 11.610 2.420 ;
        RECT  11.210 1.570 11.450 3.210 ;
        RECT  10.070 1.570 11.210 1.810 ;
        RECT  10.590 2.970 11.210 3.210 ;
        RECT  10.190 2.970 10.590 3.370 ;
        RECT  9.890 2.290 10.290 2.690 ;
        RECT  9.670 1.220 10.070 1.810 ;
        RECT  8.870 2.370 9.890 2.610 ;
        RECT  9.390 1.570 9.670 1.810 ;
        RECT  9.150 1.570 9.390 1.970 ;
        RECT  8.630 1.610 8.870 3.760 ;
        RECT  8.130 1.610 8.630 1.850 ;
        RECT  8.190 3.360 8.630 3.760 ;
        RECT  7.610 0.670 8.510 0.910 ;
        RECT  7.610 2.810 8.350 3.050 ;
        RECT  7.890 1.450 8.130 1.850 ;
        RECT  7.370 0.670 7.610 3.050 ;
        RECT  6.230 1.240 7.370 1.480 ;
        RECT  6.930 2.810 7.370 3.050 ;
        RECT  6.890 2.020 7.130 2.420 ;
        RECT  6.690 2.810 6.930 3.390 ;
        RECT  6.180 2.100 6.890 2.340 ;
        RECT  6.470 3.150 6.690 3.390 ;
        RECT  6.270 3.670 6.510 4.070 ;
        RECT  3.710 3.670 6.270 3.910 ;
        RECT  5.990 0.670 6.230 1.480 ;
        RECT  5.940 1.760 6.180 3.400 ;
        RECT  5.220 0.670 5.990 0.910 ;
        RECT  5.710 1.760 5.940 2.000 ;
        RECT  4.230 3.160 5.940 3.400 ;
        RECT  5.470 1.430 5.710 2.000 ;
        RECT  5.160 2.370 5.400 2.770 ;
        RECT  4.940 2.370 5.160 2.610 ;
        RECT  4.700 1.150 4.940 2.610 ;
        RECT  3.070 1.150 4.700 1.390 ;
        RECT  3.990 2.530 4.230 3.400 ;
        RECT  3.470 1.830 3.710 4.170 ;
        RECT  3.310 1.830 3.470 2.070 ;
        RECT  2.890 3.930 3.470 4.170 ;
        RECT  3.070 1.670 3.310 2.070 ;
        RECT  2.950 2.520 3.190 3.500 ;
        RECT  2.790 0.910 3.070 1.390 ;
        RECT  2.790 2.520 2.950 2.760 ;
        RECT  2.490 3.930 2.890 4.300 ;
        RECT  2.670 0.910 2.790 2.760 ;
        RECT  2.550 1.150 2.670 2.760 ;
        RECT  0.850 3.930 2.490 4.170 ;
        RECT  0.510 1.280 0.910 1.680 ;
        RECT  0.610 3.050 0.850 4.170 ;
        RECT  0.500 3.050 0.610 3.450 ;
        RECT  0.500 1.440 0.510 1.680 ;
        RECT  0.450 1.440 0.500 3.450 ;
        RECT  0.260 1.440 0.450 3.290 ;
    END
END DFFNSXL

MACRO DFFNSX4
    CLASS CORE ;
    FOREIGN DFFNSX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNSXL ;
    SIZE 18.480 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.070 4.060 4.690 4.380 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.290 1.260 15.330 2.660 ;
        RECT  15.330 1.260 15.730 3.200 ;
        RECT  15.730 1.260 15.760 1.660 ;
        RECT  15.730 2.800 16.140 3.200 ;
        RECT  15.760 0.660 16.160 1.660 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.200 0.860 17.240 1.260 ;
        RECT  17.260 2.800 17.270 3.200 ;
        RECT  17.240 0.860 17.270 2.180 ;
        RECT  17.270 0.860 17.600 3.220 ;
        RECT  17.600 1.820 17.710 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.450 1.820 1.870 2.520 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.760 2.010 1.170 2.660 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.920 5.440 ;
        RECT  0.920 3.710 0.930 5.440 ;
        RECT  0.930 3.590 1.330 5.440 ;
        RECT  1.330 3.710 1.340 5.440 ;
        RECT  1.340 4.640 3.560 5.440 ;
        RECT  3.560 4.170 3.800 5.440 ;
        RECT  3.800 4.640 5.010 5.440 ;
        RECT  5.010 4.310 5.020 5.440 ;
        RECT  5.020 4.190 5.420 5.440 ;
        RECT  5.420 4.310 5.430 5.440 ;
        RECT  5.430 4.640 6.350 5.440 ;
        RECT  6.350 4.030 6.360 5.440 ;
        RECT  6.360 3.830 6.760 5.440 ;
        RECT  6.760 4.030 6.770 5.440 ;
        RECT  6.770 4.640 8.870 5.440 ;
        RECT  8.870 3.630 9.270 5.440 ;
        RECT  9.270 4.640 10.720 5.440 ;
        RECT  10.720 4.010 11.120 5.440 ;
        RECT  11.120 4.640 12.230 5.440 ;
        RECT  12.230 3.490 12.630 5.440 ;
        RECT  12.630 4.640 13.670 5.440 ;
        RECT  13.670 3.490 14.070 5.440 ;
        RECT  14.070 4.640 15.110 5.440 ;
        RECT  15.110 4.010 15.510 5.440 ;
        RECT  15.510 4.640 16.500 5.440 ;
        RECT  16.500 4.210 16.510 5.440 ;
        RECT  16.510 4.010 16.910 5.440 ;
        RECT  16.910 4.210 16.920 5.440 ;
        RECT  16.920 4.640 17.900 5.440 ;
        RECT  17.900 4.210 17.910 5.440 ;
        RECT  17.910 4.010 18.310 5.440 ;
        RECT  18.310 4.210 18.320 5.440 ;
        RECT  18.320 4.640 18.480 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        RECT  0.990 -0.400 1.390 0.560 ;
        RECT  1.390 -0.400 3.590 0.400 ;
        RECT  3.590 -0.400 3.600 1.000 ;
        RECT  3.600 -0.400 4.000 1.120 ;
        RECT  4.000 -0.400 4.010 1.000 ;
        RECT  4.010 -0.400 6.490 0.400 ;
        RECT  6.490 -0.400 6.500 0.910 ;
        RECT  6.500 -0.400 6.900 1.110 ;
        RECT  6.900 -0.400 6.910 0.910 ;
        RECT  6.910 -0.400 9.120 0.400 ;
        RECT  9.120 -0.400 9.520 0.560 ;
        RECT  9.520 -0.400 11.120 0.400 ;
        RECT  11.120 -0.400 11.520 0.560 ;
        RECT  11.520 -0.400 13.600 0.400 ;
        RECT  13.600 -0.400 14.000 1.220 ;
        RECT  14.000 -0.400 15.040 0.400 ;
        RECT  15.040 -0.400 15.440 0.890 ;
        RECT  15.440 -0.400 16.480 0.400 ;
        RECT  16.480 -0.400 16.880 1.440 ;
        RECT  16.880 -0.400 17.920 0.400 ;
        RECT  17.920 -0.400 18.320 1.460 ;
        RECT  18.320 -0.400 18.480 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  17.950 2.030 18.190 3.730 ;
        RECT  15.050 3.490 17.950 3.730 ;
        RECT  14.810 1.390 15.050 3.730 ;
        RECT  14.720 1.390 14.810 1.630 ;
        RECT  14.390 2.890 14.810 3.290 ;
        RECT  14.320 1.230 14.720 1.630 ;
        RECT  13.540 2.050 14.570 2.450 ;
        RECT  13.350 1.500 13.540 3.210 ;
        RECT  13.300 1.500 13.350 3.370 ;
        RECT  12.790 1.500 13.300 1.740 ;
        RECT  12.950 2.970 13.300 3.370 ;
        RECT  12.100 2.100 13.000 2.500 ;
        RECT  11.910 2.970 12.950 3.210 ;
        RECT  12.390 1.050 12.790 1.740 ;
        RECT  10.760 1.050 12.390 1.290 ;
        RECT  10.200 2.180 12.100 2.420 ;
        RECT  11.750 2.970 11.910 3.370 ;
        RECT  11.510 2.970 11.750 3.730 ;
        RECT  10.450 3.490 11.510 3.730 ;
        RECT  10.210 3.490 10.450 4.070 ;
        RECT  8.700 0.860 10.380 1.100 ;
        RECT  10.160 1.380 10.200 2.420 ;
        RECT  9.960 1.380 10.160 3.090 ;
        RECT  9.740 1.380 9.960 1.780 ;
        RECT  9.920 2.180 9.960 3.090 ;
        RECT  9.720 2.850 9.920 3.090 ;
        RECT  8.180 1.380 9.740 1.620 ;
        RECT  9.480 2.850 9.720 3.310 ;
        RECT  9.440 2.170 9.680 2.570 ;
        RECT  8.020 3.070 9.480 3.310 ;
        RECT  8.520 2.170 9.440 2.410 ;
        RECT  8.460 0.670 8.700 1.100 ;
        RECT  8.280 1.920 8.520 2.410 ;
        RECT  7.490 0.670 8.460 0.910 ;
        RECT  8.120 1.920 8.280 2.160 ;
        RECT  7.780 1.190 8.180 1.620 ;
        RECT  7.620 3.070 8.020 3.470 ;
        RECT  7.500 2.280 7.800 2.680 ;
        RECT  7.360 2.270 7.500 2.680 ;
        RECT  7.360 0.670 7.490 1.630 ;
        RECT  7.250 0.670 7.360 3.270 ;
        RECT  7.120 1.390 7.250 3.270 ;
        RECT  6.020 1.390 7.120 1.650 ;
        RECT  5.840 3.030 7.120 3.270 ;
        RECT  5.560 2.230 6.840 2.640 ;
        RECT  5.860 1.240 6.020 1.650 ;
        RECT  5.700 3.550 5.940 4.130 ;
        RECT  5.700 0.670 5.860 1.650 ;
        RECT  5.620 0.670 5.700 1.640 ;
        RECT  3.280 3.550 5.700 3.790 ;
        RECT  5.560 0.670 5.620 1.070 ;
        RECT  5.320 1.930 5.560 3.270 ;
        RECT  5.200 1.930 5.320 2.170 ;
        RECT  3.800 3.030 5.320 3.270 ;
        RECT  4.960 0.930 5.200 2.170 ;
        RECT  4.630 2.450 5.040 2.690 ;
        RECT  4.390 1.400 4.630 2.690 ;
        RECT  2.660 1.400 4.390 1.640 ;
        RECT  3.560 2.180 3.800 3.270 ;
        RECT  3.540 2.180 3.560 2.580 ;
        RECT  3.260 2.890 3.280 4.370 ;
        RECT  3.040 1.990 3.260 4.370 ;
        RECT  3.020 1.990 3.040 3.130 ;
        RECT  1.910 4.130 3.040 4.370 ;
        RECT  2.820 1.990 3.020 2.390 ;
        RECT  2.540 3.410 2.760 3.810 ;
        RECT  2.540 0.990 2.660 1.640 ;
        RECT  2.300 0.990 2.540 3.810 ;
        RECT  2.260 0.990 2.300 1.390 ;
        RECT  1.670 2.990 1.910 4.370 ;
        RECT  0.570 2.990 1.670 3.230 ;
        RECT  0.400 1.070 0.570 1.470 ;
        RECT  0.400 2.990 0.570 3.720 ;
        RECT  0.170 1.070 0.400 3.720 ;
        RECT  0.160 1.230 0.170 3.720 ;
    END
END DFFNSX4

MACRO DFFNSX2
    CLASS CORE ;
    FOREIGN DFFNSX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNSXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.760 2.090 ;
        RECT  3.760 1.850 3.810 2.090 ;
        RECT  3.810 1.850 4.050 2.400 ;
        RECT  4.050 2.000 4.210 2.400 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.850 2.750 11.890 3.150 ;
        RECT  11.730 0.670 11.890 0.910 ;
        RECT  11.890 0.670 12.070 3.150 ;
        RECT  12.070 0.670 12.130 3.160 ;
        RECT  12.130 2.390 12.340 3.160 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.740 1.270 12.850 1.530 ;
        RECT  12.850 1.260 13.290 1.540 ;
        RECT  13.290 0.700 13.410 1.680 ;
        RECT  13.290 3.130 13.450 4.110 ;
        RECT  13.410 0.700 13.450 1.840 ;
        RECT  13.450 0.700 13.690 4.110 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.270 1.120 1.530 ;
        RECT  1.120 1.290 1.160 1.530 ;
        RECT  1.160 1.290 1.400 2.140 ;
        RECT  1.400 1.740 1.560 2.140 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.780 2.530 0.880 2.930 ;
        RECT  0.880 2.530 1.120 3.200 ;
        RECT  1.120 2.960 1.520 3.200 ;
        RECT  1.520 2.950 1.780 3.210 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.850 5.440 ;
        RECT  0.850 4.480 1.250 5.440 ;
        RECT  1.250 4.640 3.390 5.440 ;
        RECT  3.390 4.480 3.790 5.440 ;
        RECT  3.790 4.640 4.920 5.440 ;
        RECT  4.920 4.310 4.930 5.440 ;
        RECT  4.930 4.190 5.330 5.440 ;
        RECT  5.330 4.310 5.340 5.440 ;
        RECT  5.340 4.640 6.320 5.440 ;
        RECT  6.320 3.880 6.330 5.440 ;
        RECT  6.330 3.680 6.730 5.440 ;
        RECT  6.730 3.880 6.740 5.440 ;
        RECT  6.740 4.640 8.820 5.440 ;
        RECT  8.820 4.010 9.060 5.440 ;
        RECT  9.060 4.640 10.380 5.440 ;
        RECT  10.380 4.480 10.780 5.440 ;
        RECT  10.780 4.640 12.520 5.440 ;
        RECT  12.520 4.290 12.530 5.440 ;
        RECT  12.530 4.090 12.930 5.440 ;
        RECT  12.930 4.290 12.940 5.440 ;
        RECT  12.940 4.640 13.860 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.840 0.400 ;
        RECT  0.840 -0.400 1.240 0.560 ;
        RECT  1.240 -0.400 3.590 0.400 ;
        RECT  3.590 -0.400 3.600 0.910 ;
        RECT  3.600 -0.400 4.000 1.030 ;
        RECT  4.000 -0.400 4.010 0.910 ;
        RECT  4.010 -0.400 6.020 0.400 ;
        RECT  6.020 -0.400 6.260 1.110 ;
        RECT  6.260 -0.400 8.810 0.400 ;
        RECT  8.810 -0.400 9.210 1.000 ;
        RECT  9.210 -0.400 10.580 0.400 ;
        RECT  10.580 -0.400 10.980 0.560 ;
        RECT  10.980 -0.400 12.520 0.400 ;
        RECT  12.520 -0.400 12.530 0.790 ;
        RECT  12.530 -0.400 12.930 0.990 ;
        RECT  12.930 -0.400 12.940 0.790 ;
        RECT  12.940 -0.400 13.860 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  13.010 2.170 13.170 2.570 ;
        RECT  12.770 2.170 13.010 3.740 ;
        RECT  11.570 3.500 12.770 3.740 ;
        RECT  11.570 1.330 11.590 1.730 ;
        RECT  11.330 1.330 11.570 3.740 ;
        RECT  11.190 1.330 11.330 1.730 ;
        RECT  11.030 3.020 11.330 3.420 ;
        RECT  10.260 2.010 11.050 2.450 ;
        RECT  10.020 1.510 10.260 3.220 ;
        RECT  9.710 1.510 10.020 1.750 ;
        RECT  9.960 2.980 10.020 3.220 ;
        RECT  9.800 2.980 9.960 3.380 ;
        RECT  9.560 2.980 9.800 3.730 ;
        RECT  9.320 2.100 9.720 2.500 ;
        RECT  9.310 1.240 9.710 1.750 ;
        RECT  8.520 3.490 9.560 3.730 ;
        RECT  8.290 2.180 9.320 2.420 ;
        RECT  8.510 1.240 9.310 1.480 ;
        RECT  8.280 3.490 8.520 4.070 ;
        RECT  8.050 1.880 8.290 3.160 ;
        RECT  8.120 3.670 8.280 4.070 ;
        RECT  7.870 0.670 8.110 1.560 ;
        RECT  7.540 1.880 8.050 2.120 ;
        RECT  7.930 2.920 8.050 3.160 ;
        RECT  7.690 2.920 7.930 3.330 ;
        RECT  7.020 0.670 7.870 0.910 ;
        RECT  7.020 2.400 7.750 2.640 ;
        RECT  7.300 1.190 7.540 2.120 ;
        RECT  6.780 0.670 7.020 3.180 ;
        RECT  5.730 1.390 6.780 1.650 ;
        RECT  6.210 2.940 6.780 3.180 ;
        RECT  6.260 1.930 6.500 2.330 ;
        RECT  5.530 1.970 6.260 2.210 ;
        RECT  5.810 2.940 6.210 3.340 ;
        RECT  5.610 3.670 5.850 4.070 ;
        RECT  5.490 0.670 5.730 1.650 ;
        RECT  3.050 3.670 5.610 3.910 ;
        RECT  5.290 1.970 5.530 3.390 ;
        RECT  4.490 0.670 5.490 0.910 ;
        RECT  5.210 1.970 5.290 2.210 ;
        RECT  3.570 3.150 5.290 3.390 ;
        RECT  4.970 1.430 5.210 2.210 ;
        RECT  4.690 2.520 4.980 2.760 ;
        RECT  4.450 1.310 4.690 2.760 ;
        RECT  3.320 1.310 4.450 1.550 ;
        RECT  3.330 2.720 3.570 3.390 ;
        RECT  3.080 1.150 3.320 1.550 ;
        RECT  2.580 1.150 3.080 1.390 ;
        RECT  2.810 1.830 3.050 4.100 ;
        RECT  2.800 1.830 2.810 2.070 ;
        RECT  0.600 3.860 2.810 4.100 ;
        RECT  2.560 1.670 2.800 2.070 ;
        RECT  2.280 0.700 2.580 1.390 ;
        RECT  2.290 2.360 2.530 3.580 ;
        RECT  2.280 2.360 2.290 2.600 ;
        RECT  2.180 0.700 2.280 2.600 ;
        RECT  2.040 1.150 2.180 2.600 ;
        RECT  0.490 3.240 0.600 4.100 ;
        RECT  0.360 1.150 0.490 4.100 ;
        RECT  0.250 1.150 0.360 3.640 ;
        RECT  0.200 3.240 0.250 3.640 ;
    END
END DFFNSX2

MACRO DFFNSX1
    CLASS CORE ;
    FOREIGN DFFNSX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNSXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  10.010 3.930 10.570 4.350 ;
        RECT  10.570 3.940 10.640 4.340 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.700 3.650 12.000 4.050 ;
        RECT  12.000 3.510 12.100 4.050 ;
        RECT  11.700 0.670 12.100 1.100 ;
        RECT  12.100 3.500 12.240 3.890 ;
        RECT  12.240 3.500 12.340 3.770 ;
        RECT  12.340 3.500 12.660 3.740 ;
        RECT  12.100 0.860 12.660 1.100 ;
        RECT  12.660 0.860 12.900 3.740 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.290 2.840 13.310 3.240 ;
        RECT  13.290 1.220 13.310 1.620 ;
        RECT  13.310 1.210 13.700 3.250 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.440 1.280 1.450 1.760 ;
        RECT  1.450 1.280 1.520 1.840 ;
        RECT  1.520 1.270 1.850 1.840 ;
        RECT  1.850 1.270 1.860 1.770 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.830 2.290 0.950 2.690 ;
        RECT  0.950 2.280 1.280 2.700 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.480 5.440 ;
        RECT  1.480 4.480 1.880 5.440 ;
        RECT  1.880 4.640 4.220 5.440 ;
        RECT  4.220 4.480 4.620 5.440 ;
        RECT  4.620 4.640 5.640 5.440 ;
        RECT  5.640 4.210 5.650 5.440 ;
        RECT  5.650 4.090 6.050 5.440 ;
        RECT  6.050 4.210 6.060 5.440 ;
        RECT  6.060 4.640 6.950 5.440 ;
        RECT  6.950 3.790 6.960 5.440 ;
        RECT  6.960 3.590 7.360 5.440 ;
        RECT  7.360 3.790 7.370 5.440 ;
        RECT  7.370 4.640 9.290 5.440 ;
        RECT  9.290 3.790 9.300 5.440 ;
        RECT  9.300 3.590 9.700 5.440 ;
        RECT  9.700 3.790 9.710 5.440 ;
        RECT  9.710 4.640 10.910 5.440 ;
        RECT  10.880 3.080 10.910 3.480 ;
        RECT  10.910 3.070 11.330 5.440 ;
        RECT  11.330 4.640 12.490 5.440 ;
        RECT  12.490 4.480 12.890 5.440 ;
        RECT  12.890 4.640 13.860 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.150 0.400 ;
        RECT  1.150 -0.400 1.550 0.560 ;
        RECT  1.550 -0.400 3.820 0.400 ;
        RECT  3.820 -0.400 3.830 0.880 ;
        RECT  3.830 -0.400 4.230 1.000 ;
        RECT  4.230 -0.400 4.240 0.880 ;
        RECT  4.240 -0.400 6.490 0.400 ;
        RECT  6.490 -0.400 6.730 0.950 ;
        RECT  6.730 -0.400 8.870 0.400 ;
        RECT  8.870 -0.400 9.270 0.560 ;
        RECT  9.270 -0.400 10.930 0.400 ;
        RECT  10.930 -0.400 10.940 0.670 ;
        RECT  10.940 -0.400 11.340 0.870 ;
        RECT  11.340 -0.400 11.350 0.670 ;
        RECT  11.350 -0.400 12.340 0.400 ;
        RECT  12.340 -0.400 12.900 0.560 ;
        RECT  12.900 -0.400 13.860 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.140 1.380 12.380 3.230 ;
        RECT  11.760 1.380 12.140 1.780 ;
        RECT  11.760 2.990 12.140 3.230 ;
        RECT  11.180 2.110 11.580 2.510 ;
        RECT  10.520 2.190 11.180 2.430 ;
        RECT  10.280 1.630 10.520 3.430 ;
        RECT  10.060 1.630 10.280 1.870 ;
        RECT  10.120 3.030 10.280 3.430 ;
        RECT  9.660 1.160 10.060 1.870 ;
        RECT  9.760 2.350 10.000 2.750 ;
        RECT  8.500 2.510 9.760 2.750 ;
        RECT  9.220 1.630 9.660 1.870 ;
        RECT  8.820 1.630 9.220 2.030 ;
        RECT  8.500 3.520 8.580 3.920 ;
        RECT  8.260 1.350 8.500 3.920 ;
        RECT  7.470 0.670 8.450 0.910 ;
        RECT  8.150 1.350 8.260 1.590 ;
        RECT  8.180 3.520 8.260 3.920 ;
        RECT  7.750 1.190 8.150 1.590 ;
        RECT  7.470 2.510 7.980 2.920 ;
        RECT  7.230 0.670 7.470 2.920 ;
        RECT  6.170 1.230 7.230 1.470 ;
        RECT  7.030 2.680 7.230 2.920 ;
        RECT  6.630 2.680 7.030 3.180 ;
        RECT  6.310 1.750 6.950 2.150 ;
        RECT  6.410 3.570 6.650 4.070 ;
        RECT  3.930 3.570 6.410 3.810 ;
        RECT  6.070 1.750 6.310 3.290 ;
        RECT  5.930 0.670 6.170 1.470 ;
        RECT  5.650 1.750 6.070 1.990 ;
        RECT  4.470 3.050 6.070 3.290 ;
        RECT  4.510 0.670 5.930 0.910 ;
        RECT  5.390 2.370 5.790 2.770 ;
        RECT  5.410 1.370 5.650 1.990 ;
        RECT  4.990 2.370 5.390 2.610 ;
        RECT  4.750 1.280 4.990 2.610 ;
        RECT  2.890 1.280 4.750 1.520 ;
        RECT  4.230 2.130 4.470 3.290 ;
        RECT  4.170 2.130 4.230 2.370 ;
        RECT  3.930 1.970 4.170 2.370 ;
        RECT  3.690 2.650 3.930 4.090 ;
        RECT  3.190 2.650 3.690 2.890 ;
        RECT  1.050 3.850 3.690 4.090 ;
        RECT  3.170 3.160 3.410 3.560 ;
        RECT  2.950 1.800 3.190 2.890 ;
        RECT  2.510 3.160 3.170 3.400 ;
        RECT  2.790 1.800 2.950 2.040 ;
        RECT  2.510 1.000 2.890 1.520 ;
        RECT  2.490 1.000 2.510 3.400 ;
        RECT  2.270 1.280 2.490 3.400 ;
        RECT  0.810 2.970 1.050 4.090 ;
        RECT  0.650 2.970 0.810 3.370 ;
        RECT  0.500 2.970 0.650 3.210 ;
        RECT  0.500 1.330 0.570 1.730 ;
        RECT  0.260 1.330 0.500 3.210 ;
        RECT  0.170 1.330 0.260 1.730 ;
    END
END DFFNSX1

MACRO DFFNRXL
    CLASS CORE ;
    FOREIGN DFFNRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 2.390 4.290 2.650 ;
        RECT  4.290 2.390 4.420 3.190 ;
        RECT  4.420 2.400 4.530 3.190 ;
        RECT  4.530 2.940 4.730 3.190 ;
        RECT  4.730 2.950 4.970 3.190 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.320 0.720 13.330 1.100 ;
        RECT  13.190 3.690 13.590 4.090 ;
        RECT  13.330 0.710 13.730 1.100 ;
        RECT  13.590 3.690 14.120 3.930 ;
        RECT  13.730 0.860 14.120 1.100 ;
        RECT  14.120 0.860 14.360 3.930 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.690 1.380 14.720 2.070 ;
        RECT  14.690 3.040 14.730 3.460 ;
        RECT  14.720 1.380 14.730 2.090 ;
        RECT  14.730 1.380 14.930 3.460 ;
        RECT  14.930 1.830 14.970 3.460 ;
        RECT  14.970 1.830 14.980 2.090 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.460 1.510 1.900 2.090 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 0.880 2.650 ;
        RECT  0.880 2.390 1.120 2.870 ;
        RECT  1.120 2.400 1.200 2.870 ;
        RECT  1.200 2.470 1.280 2.870 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.170 5.440 ;
        RECT  1.170 4.480 1.570 5.440 ;
        RECT  1.570 4.640 4.300 5.440 ;
        RECT  4.300 4.480 4.700 5.440 ;
        RECT  4.700 4.640 7.770 5.440 ;
        RECT  7.770 4.110 8.750 5.440 ;
        RECT  8.750 4.640 11.100 5.440 ;
        RECT  11.100 4.180 11.110 5.440 ;
        RECT  11.110 3.980 11.510 5.440 ;
        RECT  11.510 4.180 11.520 5.440 ;
        RECT  11.520 4.640 14.010 5.440 ;
        RECT  14.010 4.480 14.410 5.440 ;
        RECT  14.410 4.640 15.180 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.150 0.400 ;
        RECT  1.150 -0.400 1.550 0.560 ;
        RECT  1.550 -0.400 3.970 0.400 ;
        RECT  3.970 -0.400 3.980 0.730 ;
        RECT  3.980 -0.400 4.380 0.850 ;
        RECT  4.380 -0.400 4.390 0.730 ;
        RECT  4.390 -0.400 6.070 0.400 ;
        RECT  6.070 -0.400 6.380 1.540 ;
        RECT  6.380 1.190 6.630 1.530 ;
        RECT  6.630 1.190 7.880 1.540 ;
        RECT  7.880 1.190 8.280 1.880 ;
        RECT  6.380 -0.400 10.560 0.400 ;
        RECT  10.560 -0.400 10.570 1.110 ;
        RECT  10.570 -0.400 10.970 1.310 ;
        RECT  10.970 -0.400 10.980 1.110 ;
        RECT  10.980 -0.400 12.440 0.400 ;
        RECT  12.440 -0.400 12.450 0.690 ;
        RECT  12.450 -0.400 12.850 0.890 ;
        RECT  12.850 -0.400 12.860 0.690 ;
        RECT  12.860 -0.400 14.410 0.400 ;
        RECT  14.410 -0.400 14.810 0.560 ;
        RECT  14.810 -0.400 15.180 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  13.600 1.450 13.840 3.150 ;
        RECT  13.330 1.450 13.600 1.690 ;
        RECT  13.450 2.910 13.600 3.150 ;
        RECT  13.210 2.910 13.450 3.340 ;
        RECT  12.900 1.970 13.200 2.370 ;
        RECT  12.790 1.590 12.900 3.590 ;
        RECT  12.660 1.590 12.790 3.750 ;
        RECT  11.970 1.590 12.660 1.830 ;
        RECT  12.390 3.350 12.660 3.750 ;
        RECT  11.980 2.110 12.380 2.510 ;
        RECT  10.550 2.270 11.980 2.510 ;
        RECT  11.570 1.130 11.970 1.830 ;
        RECT  10.670 1.590 11.570 1.830 ;
        RECT  10.270 1.590 10.670 1.940 ;
        RECT  10.310 2.270 10.550 3.780 ;
        RECT  9.480 2.270 10.310 2.510 ;
        RECT  10.290 3.540 10.310 3.780 ;
        RECT  9.890 3.540 10.290 3.940 ;
        RECT  9.630 2.790 10.030 3.100 ;
        RECT  8.940 0.670 9.920 0.910 ;
        RECT  8.940 2.790 9.630 3.030 ;
        RECT  9.240 1.330 9.480 2.510 ;
        RECT  8.700 0.670 8.940 3.030 ;
        RECT  6.650 0.670 8.700 0.910 ;
        RECT  8.460 2.760 8.700 3.030 ;
        RECT  8.220 2.760 8.460 3.450 ;
        RECT  6.890 2.230 8.420 2.470 ;
        RECT  7.650 2.870 7.890 3.830 ;
        RECT  7.500 3.590 7.650 3.830 ;
        RECT  7.260 3.590 7.500 4.370 ;
        RECT  5.210 4.130 7.260 4.370 ;
        RECT  6.650 1.820 6.890 3.690 ;
        RECT  5.800 1.820 6.650 2.060 ;
        RECT  6.550 3.450 6.650 3.690 ;
        RECT  6.150 3.450 6.550 3.850 ;
        RECT  5.730 2.340 6.370 2.580 ;
        RECT  5.560 1.110 5.800 2.060 ;
        RECT  5.490 2.340 5.730 3.850 ;
        RECT  5.430 1.110 5.560 1.890 ;
        RECT  5.280 2.340 5.490 2.580 ;
        RECT  3.930 1.650 5.430 1.890 ;
        RECT  4.880 2.170 5.280 2.580 ;
        RECT  4.970 3.940 5.210 4.370 ;
        RECT  4.900 0.770 5.130 1.010 ;
        RECT  3.800 3.940 4.970 4.180 ;
        RECT  4.660 0.770 4.900 1.370 ;
        RECT  2.890 1.130 4.660 1.370 ;
        RECT  3.530 1.650 3.930 2.110 ;
        RECT  3.560 2.390 3.800 4.180 ;
        RECT  3.250 2.390 3.560 2.630 ;
        RECT  2.910 3.940 3.560 4.180 ;
        RECT  3.010 1.710 3.250 2.630 ;
        RECT  2.610 3.420 3.150 3.660 ;
        RECT  2.890 1.710 3.010 2.110 ;
        RECT  2.510 3.940 2.910 4.370 ;
        RECT  2.610 0.950 2.890 1.370 ;
        RECT  2.370 0.950 2.610 3.660 ;
        RECT  0.590 3.940 2.510 4.180 ;
        RECT  0.500 1.270 0.590 1.670 ;
        RECT  0.500 3.170 0.590 4.180 ;
        RECT  0.350 1.270 0.500 4.180 ;
        RECT  0.260 1.270 0.350 3.570 ;
        RECT  0.190 1.270 0.260 1.670 ;
        RECT  0.190 3.170 0.260 3.570 ;
    END
END DFFNRXL

MACRO DFFNRX4
    CLASS CORE ;
    FOREIGN DFFNRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNRXL ;
    SIZE 19.800 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.040 2.810 4.510 3.220 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  17.170 1.170 17.250 1.570 ;
        RECT  16.990 2.750 17.270 3.150 ;
        RECT  17.250 1.170 17.270 2.070 ;
        RECT  17.270 1.170 17.490 3.220 ;
        RECT  17.490 1.170 17.570 1.570 ;
        RECT  17.490 1.820 17.710 3.220 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  18.510 2.750 18.540 3.150 ;
        RECT  18.540 2.610 18.590 3.150 ;
        RECT  18.520 1.170 18.590 1.570 ;
        RECT  18.590 1.170 18.910 3.150 ;
        RECT  18.910 1.170 18.920 3.070 ;
        RECT  18.920 1.250 18.930 3.070 ;
        RECT  18.930 1.260 19.030 2.660 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.310 2.380 1.870 2.720 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.670 2.000 0.680 2.420 ;
        RECT  0.680 1.840 0.860 2.420 ;
        RECT  0.860 1.830 0.930 2.420 ;
        RECT  0.930 1.830 1.120 2.090 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.940 5.440 ;
        RECT  0.940 4.480 1.340 5.440 ;
        RECT  1.340 4.640 3.500 5.440 ;
        RECT  3.500 4.480 3.900 5.440 ;
        RECT  3.900 4.640 7.120 5.440 ;
        RECT  7.120 3.910 7.130 5.440 ;
        RECT  7.130 3.710 7.530 5.440 ;
        RECT  7.530 3.910 7.540 5.440 ;
        RECT  7.540 4.640 9.850 5.440 ;
        RECT  9.850 3.730 10.250 5.440 ;
        RECT  10.250 4.640 12.520 5.440 ;
        RECT  12.520 4.170 12.920 5.440 ;
        RECT  12.920 4.640 14.940 5.440 ;
        RECT  14.940 3.090 15.340 5.440 ;
        RECT  15.340 4.640 16.380 5.440 ;
        RECT  16.380 4.010 16.780 5.440 ;
        RECT  16.780 4.640 17.830 5.440 ;
        RECT  17.830 4.210 17.840 5.440 ;
        RECT  17.840 4.010 18.240 5.440 ;
        RECT  18.240 4.210 18.250 5.440 ;
        RECT  18.250 4.640 19.180 5.440 ;
        RECT  19.180 4.010 19.580 5.440 ;
        RECT  19.580 4.640 19.800 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        RECT  0.990 -0.400 1.390 0.560 ;
        RECT  1.390 -0.400 4.370 0.400 ;
        RECT  4.370 -0.400 5.350 1.290 ;
        RECT  5.350 -0.400 6.290 0.400 ;
        RECT  6.290 -0.400 6.300 0.890 ;
        RECT  6.300 -0.400 6.700 1.090 ;
        RECT  6.700 -0.400 6.710 0.890 ;
        RECT  6.710 -0.400 7.990 0.400 ;
        RECT  7.990 -0.400 8.000 1.110 ;
        RECT  8.000 -0.400 8.400 1.310 ;
        RECT  8.400 -0.400 8.410 1.110 ;
        RECT  8.410 -0.400 10.900 0.400 ;
        RECT  10.900 -0.400 11.300 0.560 ;
        RECT  11.300 -0.400 12.290 0.400 ;
        RECT  12.290 -0.400 12.300 0.710 ;
        RECT  12.300 -0.400 12.700 0.910 ;
        RECT  12.700 -0.400 12.710 0.710 ;
        RECT  12.710 -0.400 13.760 0.400 ;
        RECT  13.760 -0.400 14.160 0.910 ;
        RECT  14.160 -0.400 15.200 0.400 ;
        RECT  15.200 -0.400 15.600 0.910 ;
        RECT  15.600 -0.400 16.550 0.400 ;
        RECT  16.550 -0.400 16.560 0.690 ;
        RECT  16.560 -0.400 16.960 0.890 ;
        RECT  16.960 -0.400 16.970 0.690 ;
        RECT  16.970 -0.400 17.830 0.400 ;
        RECT  17.830 -0.400 17.840 0.690 ;
        RECT  17.840 -0.400 18.240 0.890 ;
        RECT  18.240 -0.400 18.250 0.690 ;
        RECT  18.250 -0.400 19.190 0.400 ;
        RECT  19.190 -0.400 19.590 0.890 ;
        RECT  19.590 -0.400 19.800 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  19.270 2.180 19.510 3.730 ;
        RECT  16.750 3.490 19.270 3.730 ;
        RECT  16.510 1.550 16.750 3.730 ;
        RECT  16.320 1.550 16.510 1.790 ;
        RECT  16.060 3.020 16.510 3.730 ;
        RECT  15.920 1.390 16.320 1.790 ;
        RECT  15.290 2.070 16.270 2.470 ;
        RECT  15.660 3.020 16.060 4.000 ;
        RECT  14.840 2.150 15.290 2.390 ;
        RECT  14.840 0.690 14.880 1.090 ;
        RECT  14.700 0.690 14.840 2.640 ;
        RECT  14.600 0.690 14.700 3.200 ;
        RECT  14.480 0.690 14.600 1.480 ;
        RECT  14.460 2.400 14.600 3.200 ;
        RECT  13.440 1.240 14.480 1.480 ;
        RECT  14.160 2.960 14.460 3.200 ;
        RECT  13.380 1.760 14.360 2.160 ;
        RECT  13.760 2.960 14.160 3.940 ;
        RECT  12.230 3.650 13.760 3.890 ;
        RECT  13.200 0.670 13.440 1.480 ;
        RECT  12.470 1.870 13.380 2.110 ;
        RECT  13.040 0.670 13.200 1.070 ;
        RECT  12.320 1.550 12.470 2.110 ;
        RECT  12.080 1.380 12.320 3.370 ;
        RECT  11.990 3.650 12.230 4.350 ;
        RECT  11.110 1.380 12.080 1.790 ;
        RECT  11.500 3.130 12.080 3.370 ;
        RECT  10.620 0.860 11.870 1.100 ;
        RECT  11.270 2.450 11.670 2.850 ;
        RECT  11.140 3.130 11.500 4.230 ;
        RECT  9.580 2.450 11.270 2.690 ;
        RECT  9.590 3.130 11.140 3.370 ;
        RECT  11.100 3.830 11.140 4.230 ;
        RECT  10.100 1.380 11.110 1.620 ;
        RECT  10.380 0.700 10.620 1.100 ;
        RECT  8.940 0.700 10.380 0.940 ;
        RECT  9.810 1.220 10.100 1.620 ;
        RECT  9.220 1.220 9.810 1.460 ;
        RECT  9.350 3.130 9.590 3.860 ;
        RECT  9.340 1.750 9.580 2.690 ;
        RECT  9.070 3.620 9.350 3.860 ;
        RECT  8.670 3.620 9.070 4.020 ;
        RECT  8.940 1.750 9.020 3.140 ;
        RECT  8.780 0.700 8.940 3.140 ;
        RECT  8.700 0.700 8.780 1.990 ;
        RECT  8.450 2.900 8.780 3.140 ;
        RECT  7.440 1.750 8.700 1.990 ;
        RECT  6.880 2.270 8.540 2.510 ;
        RECT  8.350 2.900 8.450 3.340 ;
        RECT  8.210 2.900 8.350 4.130 ;
        RECT  8.110 3.100 8.210 4.130 ;
        RECT  7.950 3.730 8.110 4.130 ;
        RECT  7.330 2.810 7.730 3.430 ;
        RECT  7.200 0.670 7.440 1.990 ;
        RECT  6.850 3.190 7.330 3.430 ;
        RECT  6.980 0.670 7.200 0.910 ;
        RECT  6.640 1.570 6.880 2.910 ;
        RECT  6.610 3.190 6.850 4.370 ;
        RECT  4.060 1.570 6.640 1.810 ;
        RECT  6.230 2.670 6.640 2.910 ;
        RECT  4.420 4.130 6.610 4.370 ;
        RECT  5.100 2.150 6.360 2.390 ;
        RECT  5.990 2.670 6.230 3.800 ;
        RECT  5.830 3.560 5.990 3.800 ;
        RECT  4.860 2.090 5.100 3.850 ;
        RECT  4.340 2.090 4.860 2.330 ;
        RECT  4.700 3.610 4.860 3.850 ;
        RECT  4.180 3.940 4.420 4.370 ;
        RECT  3.170 3.940 4.180 4.180 ;
        RECT  3.820 0.690 4.060 1.290 ;
        RECT  3.820 1.570 4.060 2.530 ;
        RECT  2.660 1.050 3.820 1.290 ;
        RECT  3.620 2.290 3.820 2.530 ;
        RECT  3.380 2.290 3.620 2.690 ;
        RECT  2.930 3.010 3.170 4.290 ;
        RECT  2.900 3.010 2.930 3.250 ;
        RECT  2.410 4.050 2.930 4.290 ;
        RECT  2.660 1.840 2.900 3.250 ;
        RECT  2.420 1.050 2.660 1.560 ;
        RECT  2.380 3.530 2.650 3.770 ;
        RECT  2.380 1.320 2.420 1.560 ;
        RECT  2.010 4.050 2.410 4.340 ;
        RECT  2.140 1.320 2.380 3.770 ;
        RECT  1.860 4.050 2.010 4.290 ;
        RECT  1.620 3.300 1.860 4.290 ;
        RECT  0.570 3.300 1.620 3.540 ;
        RECT  0.400 1.150 0.570 1.550 ;
        RECT  0.400 3.140 0.570 3.540 ;
        RECT  0.160 1.150 0.400 3.540 ;
    END
END DFFNRX4

MACRO DFFNRX2
    CLASS CORE ;
    FOREIGN DFFNRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNRXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 2.950 4.170 3.210 ;
        RECT  4.170 2.710 4.420 3.210 ;
        RECT  4.420 2.710 4.920 3.110 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.400 2.920 14.480 3.320 ;
        RECT  14.480 2.610 14.490 3.320 ;
        RECT  14.400 0.730 14.490 1.710 ;
        RECT  14.490 0.730 14.730 3.320 ;
        RECT  14.730 2.390 14.800 3.320 ;
        RECT  14.730 0.730 14.800 1.710 ;
        RECT  14.800 2.390 14.980 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.930 0.730 16.040 1.960 ;
        RECT  15.930 3.170 16.050 4.150 ;
        RECT  16.040 0.730 16.050 2.090 ;
        RECT  16.050 0.730 16.290 4.150 ;
        RECT  16.290 0.730 16.300 2.090 ;
        RECT  16.290 3.170 16.330 4.150 ;
        RECT  16.300 0.730 16.330 1.960 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.480 1.140 1.780 1.840 ;
        RECT  1.780 1.140 1.880 1.830 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.840 1.840 0.860 2.640 ;
        RECT  0.860 1.830 1.080 2.640 ;
        RECT  1.080 1.830 1.120 2.090 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.200 5.440 ;
        RECT  1.200 4.480 1.600 5.440 ;
        RECT  1.600 4.640 4.010 5.440 ;
        RECT  4.010 4.480 4.410 5.440 ;
        RECT  4.410 4.640 7.310 5.440 ;
        RECT  7.310 4.010 8.850 5.440 ;
        RECT  8.850 4.640 10.870 5.440 ;
        RECT  10.870 4.110 10.880 5.440 ;
        RECT  10.880 3.910 11.280 5.440 ;
        RECT  11.280 4.110 11.290 5.440 ;
        RECT  11.290 4.640 12.830 5.440 ;
        RECT  12.830 3.500 12.840 5.440 ;
        RECT  12.840 3.300 13.240 5.440 ;
        RECT  13.240 3.500 13.250 5.440 ;
        RECT  13.250 4.640 15.160 5.440 ;
        RECT  15.160 4.320 15.170 5.440 ;
        RECT  15.170 4.120 15.570 5.440 ;
        RECT  15.570 4.320 15.580 5.440 ;
        RECT  15.580 4.640 16.500 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.140 0.400 ;
        RECT  1.140 -0.400 1.540 0.560 ;
        RECT  1.540 -0.400 4.870 0.400 ;
        RECT  4.870 -0.400 5.270 1.310 ;
        RECT  5.270 -0.400 6.360 0.400 ;
        RECT  6.360 -0.400 6.370 0.640 ;
        RECT  6.370 -0.400 6.770 0.930 ;
        RECT  6.770 -0.400 6.780 0.640 ;
        RECT  6.780 -0.400 8.060 0.400 ;
        RECT  8.060 -0.400 8.070 1.020 ;
        RECT  8.070 -0.400 8.470 1.140 ;
        RECT  8.470 -0.400 8.480 1.020 ;
        RECT  8.480 -0.400 11.150 0.400 ;
        RECT  11.150 -0.400 11.550 0.560 ;
        RECT  11.550 -0.400 12.720 0.400 ;
        RECT  12.720 -0.400 12.730 1.100 ;
        RECT  12.730 -0.400 13.130 1.300 ;
        RECT  13.130 -0.400 13.140 1.100 ;
        RECT  13.140 -0.400 15.160 0.400 ;
        RECT  15.160 -0.400 15.170 1.200 ;
        RECT  15.170 -0.400 15.570 1.690 ;
        RECT  15.570 -0.400 15.580 1.200 ;
        RECT  15.580 -0.400 16.500 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  15.650 2.200 15.680 2.600 ;
        RECT  15.410 2.200 15.650 3.840 ;
        RECT  14.120 3.600 15.410 3.840 ;
        RECT  13.880 1.080 14.120 3.840 ;
        RECT  13.550 1.080 13.880 1.480 ;
        RECT  13.660 2.920 13.880 3.320 ;
        RECT  12.650 1.950 13.640 2.350 ;
        RECT  12.410 1.580 12.650 3.020 ;
        RECT  12.370 1.580 12.410 1.820 ;
        RECT  12.020 2.780 12.410 3.020 ;
        RECT  11.970 0.940 12.370 1.820 ;
        RECT  11.730 2.100 12.130 2.500 ;
        RECT  11.620 2.780 12.020 3.900 ;
        RECT  11.100 1.580 11.970 1.820 ;
        RECT  10.420 2.260 11.730 2.500 ;
        RECT  10.780 2.780 11.620 3.020 ;
        RECT  10.700 1.580 11.100 1.980 ;
        RECT  10.180 2.090 10.420 3.490 ;
        RECT  9.670 2.090 10.180 2.330 ;
        RECT  10.140 3.250 10.180 3.490 ;
        RECT  9.740 3.250 10.140 3.650 ;
        RECT  9.120 0.670 10.080 0.910 ;
        RECT  9.200 2.610 9.900 2.850 ;
        RECT  9.430 1.230 9.670 2.330 ;
        RECT  9.120 2.610 9.200 3.270 ;
        RECT  8.880 0.670 9.120 3.270 ;
        RECT  7.590 1.420 8.880 1.710 ;
        RECT  8.300 3.030 8.880 3.270 ;
        RECT  8.400 1.990 8.640 2.390 ;
        RECT  6.850 1.990 8.400 2.230 ;
        RECT  7.900 3.030 8.300 3.430 ;
        RECT  7.380 2.510 7.960 2.750 ;
        RECT  7.460 1.310 7.590 1.710 ;
        RECT  7.450 0.880 7.460 1.710 ;
        RECT  7.190 0.670 7.450 1.710 ;
        RECT  7.140 2.510 7.380 3.730 ;
        RECT  7.050 0.670 7.190 0.910 ;
        RECT  6.940 3.490 7.140 3.730 ;
        RECT  6.700 3.490 6.940 4.310 ;
        RECT  6.610 1.590 6.850 3.190 ;
        RECT  4.930 4.070 6.700 4.310 ;
        RECT  6.190 1.590 6.610 1.830 ;
        RECT  6.380 2.950 6.610 3.190 ;
        RECT  6.140 2.950 6.380 3.790 ;
        RECT  6.090 2.110 6.330 2.510 ;
        RECT  5.790 1.270 6.190 1.830 ;
        RECT  5.980 3.390 6.140 3.790 ;
        RECT  5.450 2.110 6.090 2.350 ;
        RECT  3.930 1.590 5.790 1.830 ;
        RECT  5.210 2.110 5.450 3.790 ;
        RECT  4.910 2.110 5.210 2.350 ;
        RECT  4.690 3.940 4.930 4.310 ;
        RECT  3.710 3.940 4.690 4.180 ;
        RECT  4.190 0.690 4.590 1.200 ;
        RECT  2.890 0.960 4.190 1.200 ;
        RECT  3.690 1.590 3.930 2.270 ;
        RECT  3.470 2.560 3.710 4.250 ;
        RECT  3.530 1.870 3.690 2.270 ;
        RECT  3.250 2.560 3.470 2.800 ;
        RECT  2.190 4.010 3.470 4.250 ;
        RECT  3.010 1.480 3.250 2.800 ;
        RECT  2.950 3.090 3.190 3.490 ;
        RECT  2.890 1.480 3.010 1.880 ;
        RECT  2.730 3.090 2.950 3.330 ;
        RECT  2.600 0.800 2.890 1.200 ;
        RECT  2.600 2.160 2.730 3.330 ;
        RECT  2.490 0.800 2.600 3.330 ;
        RECT  2.360 0.800 2.490 2.400 ;
        RECT  1.950 3.080 2.190 4.250 ;
        RECT  0.790 3.080 1.950 3.320 ;
        RECT  0.500 2.920 0.790 3.320 ;
        RECT  0.490 0.960 0.500 3.320 ;
        RECT  0.260 0.880 0.490 3.320 ;
        RECT  0.250 0.880 0.260 1.280 ;
    END
END DFFNRX2

MACRO DFFNRX1
    CLASS CORE ;
    FOREIGN DFFNRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNRXL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 2.390 4.290 2.650 ;
        RECT  4.290 2.390 4.420 3.190 ;
        RECT  4.420 2.400 4.530 3.190 ;
        RECT  4.530 2.940 4.730 3.190 ;
        RECT  4.730 2.950 4.970 3.190 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.190 3.690 13.590 4.090 ;
        RECT  13.210 0.710 13.660 1.100 ;
        RECT  13.590 3.690 14.120 3.930 ;
        RECT  13.660 0.860 14.120 1.100 ;
        RECT  14.120 0.860 14.360 3.930 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.690 1.310 14.720 2.070 ;
        RECT  14.690 3.170 14.730 3.570 ;
        RECT  14.720 1.310 14.730 2.090 ;
        RECT  14.730 1.310 14.930 3.570 ;
        RECT  14.930 1.830 14.970 3.570 ;
        RECT  14.970 1.830 14.980 2.090 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.450 1.740 1.930 2.330 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 0.870 3.210 ;
        RECT  0.870 2.640 1.120 3.210 ;
        RECT  1.120 2.640 1.410 3.040 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.470 5.440 ;
        RECT  1.470 4.480 1.870 5.440 ;
        RECT  1.870 4.640 4.290 5.440 ;
        RECT  4.290 4.480 4.690 5.440 ;
        RECT  4.690 4.640 7.770 5.440 ;
        RECT  7.770 4.110 8.750 5.440 ;
        RECT  8.750 4.640 10.690 5.440 ;
        RECT  10.690 4.190 10.700 5.440 ;
        RECT  10.700 3.990 11.100 5.440 ;
        RECT  11.100 4.190 11.110 5.440 ;
        RECT  11.110 4.640 14.010 5.440 ;
        RECT  14.010 4.480 14.410 5.440 ;
        RECT  14.410 4.640 15.180 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.160 0.400 ;
        RECT  1.160 -0.400 1.560 0.560 ;
        RECT  1.560 -0.400 3.970 0.400 ;
        RECT  3.970 -0.400 3.980 0.730 ;
        RECT  3.980 -0.400 4.380 0.850 ;
        RECT  4.380 -0.400 4.390 0.730 ;
        RECT  4.390 -0.400 6.130 0.400 ;
        RECT  6.130 -0.400 6.370 1.530 ;
        RECT  6.370 1.190 6.630 1.530 ;
        RECT  6.630 1.190 7.880 1.540 ;
        RECT  7.880 1.190 8.280 1.880 ;
        RECT  6.370 -0.400 10.560 0.400 ;
        RECT  10.560 -0.400 10.570 1.110 ;
        RECT  10.570 -0.400 10.970 1.310 ;
        RECT  10.970 -0.400 10.980 1.110 ;
        RECT  10.980 -0.400 12.440 0.400 ;
        RECT  12.440 -0.400 12.450 0.690 ;
        RECT  12.450 -0.400 12.850 0.890 ;
        RECT  12.850 -0.400 12.860 0.690 ;
        RECT  12.860 -0.400 14.500 0.400 ;
        RECT  14.500 -0.400 14.900 0.560 ;
        RECT  14.900 -0.400 15.180 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  13.600 1.450 13.840 3.150 ;
        RECT  13.270 1.450 13.600 1.690 ;
        RECT  13.450 2.910 13.600 3.150 ;
        RECT  13.210 2.910 13.450 3.340 ;
        RECT  12.900 1.970 13.200 2.370 ;
        RECT  12.780 1.590 12.900 3.590 ;
        RECT  12.660 1.590 12.780 3.750 ;
        RECT  11.970 1.590 12.660 1.830 ;
        RECT  12.380 3.350 12.660 3.750 ;
        RECT  11.980 2.110 12.380 2.510 ;
        RECT  10.290 2.270 11.980 2.510 ;
        RECT  11.570 1.020 11.970 1.830 ;
        RECT  10.950 1.590 11.570 1.830 ;
        RECT  10.550 1.590 10.950 1.990 ;
        RECT  10.230 2.270 10.290 4.130 ;
        RECT  9.990 1.420 10.230 4.130 ;
        RECT  9.540 1.420 9.990 1.660 ;
        RECT  9.890 3.730 9.990 4.130 ;
        RECT  8.940 0.670 9.920 0.910 ;
        RECT  9.460 2.470 9.700 3.000 ;
        RECT  9.300 1.260 9.540 1.660 ;
        RECT  8.940 2.760 9.460 3.000 ;
        RECT  8.700 0.670 8.940 3.000 ;
        RECT  6.650 0.670 8.700 0.910 ;
        RECT  8.460 2.760 8.700 3.000 ;
        RECT  8.220 2.760 8.460 3.450 ;
        RECT  6.980 2.230 8.420 2.470 ;
        RECT  7.650 2.870 7.890 3.830 ;
        RECT  7.500 3.590 7.650 3.830 ;
        RECT  7.260 3.590 7.500 4.370 ;
        RECT  5.210 4.130 7.260 4.370 ;
        RECT  6.740 1.820 6.980 3.390 ;
        RECT  5.850 1.820 6.740 2.060 ;
        RECT  6.470 3.150 6.740 3.390 ;
        RECT  6.230 3.150 6.470 3.850 ;
        RECT  5.730 2.340 6.460 2.580 ;
        RECT  5.610 1.110 5.850 2.060 ;
        RECT  5.490 2.340 5.730 3.850 ;
        RECT  5.430 1.110 5.610 1.890 ;
        RECT  5.280 2.340 5.490 2.580 ;
        RECT  3.930 1.650 5.430 1.890 ;
        RECT  4.880 2.170 5.280 2.580 ;
        RECT  4.970 3.940 5.210 4.370 ;
        RECT  4.900 0.770 5.130 1.010 ;
        RECT  4.010 3.940 4.970 4.180 ;
        RECT  4.660 0.770 4.900 1.370 ;
        RECT  2.890 1.130 4.660 1.370 ;
        RECT  3.800 2.930 4.010 4.360 ;
        RECT  3.530 1.650 3.930 2.110 ;
        RECT  3.770 2.390 3.800 4.360 ;
        RECT  3.560 2.390 3.770 3.170 ;
        RECT  2.620 4.120 3.770 4.360 ;
        RECT  3.120 2.390 3.560 2.630 ;
        RECT  3.220 3.510 3.490 3.750 ;
        RECT  2.980 3.420 3.220 3.750 ;
        RECT  2.880 1.980 3.120 2.630 ;
        RECT  2.600 3.420 2.980 3.660 ;
        RECT  2.600 1.130 2.890 1.700 ;
        RECT  2.380 3.940 2.620 4.360 ;
        RECT  2.380 1.130 2.600 3.660 ;
        RECT  2.360 1.460 2.380 3.660 ;
        RECT  1.030 3.940 2.380 4.180 ;
        RECT  0.790 3.490 1.030 4.180 ;
        RECT  0.630 3.490 0.790 3.890 ;
        RECT  0.500 3.490 0.630 3.730 ;
        RECT  0.500 1.360 0.580 1.760 ;
        RECT  0.260 1.360 0.500 3.730 ;
        RECT  0.180 1.360 0.260 1.760 ;
    END
END DFFNRX1

MACRO DFFNXL
    CLASS CORE ;
    FOREIGN DFFNXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  10.670 1.780 10.680 3.250 ;
        RECT  10.680 1.390 11.010 3.250 ;
        RECT  11.010 1.780 11.020 3.250 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.090 2.920 9.490 3.320 ;
        RECT  9.490 2.950 9.700 3.210 ;
        RECT  9.480 0.720 9.880 1.100 ;
        RECT  9.700 2.950 10.160 3.190 ;
        RECT  9.880 0.860 10.160 1.100 ;
        RECT  10.160 0.860 10.400 3.190 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.350 1.850 1.520 2.480 ;
        RECT  1.520 1.830 1.590 2.480 ;
        RECT  1.590 1.830 1.780 2.090 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.800 1.210 3.220 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.090 5.440 ;
        RECT  1.090 4.480 1.490 5.440 ;
        RECT  1.490 4.640 5.830 5.440 ;
        RECT  5.830 4.480 6.230 5.440 ;
        RECT  6.230 4.640 8.270 5.440 ;
        RECT  8.270 4.480 8.670 5.440 ;
        RECT  8.670 4.640 9.880 5.440 ;
        RECT  9.880 4.480 10.280 5.440 ;
        RECT  10.280 4.640 11.220 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.960 0.400 ;
        RECT  0.960 -0.400 1.360 0.560 ;
        RECT  1.360 -0.400 3.490 0.400 ;
        RECT  3.490 -0.400 3.500 0.850 ;
        RECT  3.500 -0.400 3.900 0.970 ;
        RECT  3.900 -0.400 3.910 0.850 ;
        RECT  3.910 -0.400 5.990 0.400 ;
        RECT  5.990 -0.400 6.000 1.380 ;
        RECT  6.000 -0.400 6.400 1.500 ;
        RECT  6.400 -0.400 6.410 1.380 ;
        RECT  6.410 -0.400 8.590 0.400 ;
        RECT  8.590 -0.400 8.600 0.880 ;
        RECT  8.600 -0.400 9.000 1.080 ;
        RECT  9.000 -0.400 9.010 0.880 ;
        RECT  9.010 -0.400 10.430 0.400 ;
        RECT  10.430 -0.400 10.830 0.560 ;
        RECT  10.830 -0.400 11.220 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  9.640 1.460 9.880 2.640 ;
        RECT  9.480 1.460 9.640 1.700 ;
        RECT  8.440 2.400 9.640 2.640 ;
        RECT  9.150 3.800 9.550 4.200 ;
        RECT  9.080 1.870 9.240 2.110 ;
        RECT  8.400 3.800 9.150 4.040 ;
        RECT  8.840 1.610 9.080 2.110 ;
        RECT  7.720 1.610 8.840 1.850 ;
        RECT  8.400 2.310 8.440 2.710 ;
        RECT  8.160 2.310 8.400 4.040 ;
        RECT  8.040 2.310 8.160 2.710 ;
        RECT  6.940 0.710 7.950 0.950 ;
        RECT  7.620 1.440 7.720 4.220 ;
        RECT  7.480 1.280 7.620 4.220 ;
        RECT  7.220 1.280 7.480 1.680 ;
        RECT  7.170 3.820 7.480 4.220 ;
        RECT  6.940 2.610 7.170 3.010 ;
        RECT  6.890 0.710 6.940 3.010 ;
        RECT  6.700 0.710 6.890 4.180 ;
        RECT  5.520 1.800 6.700 2.040 ;
        RECT  6.650 2.770 6.700 4.180 ;
        RECT  5.550 3.940 6.650 4.180 ;
        RECT  6.130 2.320 6.370 3.660 ;
        RECT  5.030 3.420 6.130 3.660 ;
        RECT  5.310 3.940 5.550 4.370 ;
        RECT  5.350 1.170 5.520 2.040 ;
        RECT  5.120 1.170 5.350 3.140 ;
        RECT  3.220 4.130 5.310 4.370 ;
        RECT  5.110 1.250 5.120 3.140 ;
        RECT  4.830 3.420 5.030 3.850 ;
        RECT  4.590 1.250 4.830 3.850 ;
        RECT  4.380 1.250 4.590 1.650 ;
        RECT  3.640 2.620 4.590 2.860 ;
        RECT  4.070 1.930 4.310 2.330 ;
        RECT  2.910 1.930 4.070 2.170 ;
        RECT  3.240 2.460 3.640 2.860 ;
        RECT  2.820 3.970 3.220 4.370 ;
        RECT  2.820 1.450 2.910 3.340 ;
        RECT  1.920 0.680 2.860 0.920 ;
        RECT  2.670 1.450 2.820 3.420 ;
        RECT  2.300 3.970 2.820 4.210 ;
        RECT  2.600 1.450 2.670 1.690 ;
        RECT  2.580 3.020 2.670 3.420 ;
        RECT  2.200 1.290 2.600 1.690 ;
        RECT  2.300 2.020 2.380 2.740 ;
        RECT  2.140 2.020 2.300 4.210 ;
        RECT  2.060 2.500 2.140 4.210 ;
        RECT  1.680 0.680 1.920 1.530 ;
        RECT  0.570 1.290 1.680 1.530 ;
        RECT  0.400 1.290 0.570 1.690 ;
        RECT  0.400 3.560 0.570 3.800 ;
        RECT  0.160 1.290 0.400 3.800 ;
    END
END DFFNXL

MACRO DFFNX4
    CLASS CORE ;
    FOREIGN DFFNX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNXL ;
    SIZE 16.500 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.630 1.820 15.020 3.220 ;
        RECT  15.020 1.410 15.030 3.220 ;
        RECT  15.030 1.210 15.430 3.270 ;
        RECT  15.430 1.410 15.440 3.070 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.310 1.820 13.480 3.220 ;
        RECT  13.480 1.410 13.490 3.220 ;
        RECT  13.490 1.210 13.890 3.270 ;
        RECT  13.890 1.410 13.900 3.070 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 0.880 3.210 ;
        RECT  0.880 2.940 1.120 3.210 ;
        RECT  1.120 2.940 1.450 3.180 ;
        RECT  1.450 2.370 1.690 3.180 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.690 1.840 0.930 2.280 ;
        RECT  0.930 1.840 1.520 2.080 ;
        RECT  1.520 1.830 1.780 2.090 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.030 5.440 ;
        RECT  1.030 4.480 1.430 5.440 ;
        RECT  1.430 4.640 3.630 5.440 ;
        RECT  3.630 4.480 4.030 5.440 ;
        RECT  4.030 4.640 6.180 5.440 ;
        RECT  6.180 4.480 6.580 5.440 ;
        RECT  6.580 4.640 8.680 5.440 ;
        RECT  8.680 4.140 9.080 5.440 ;
        RECT  9.080 4.640 11.270 5.440 ;
        RECT  11.270 4.480 11.670 5.440 ;
        RECT  11.670 4.640 12.870 5.440 ;
        RECT  12.870 4.270 12.880 5.440 ;
        RECT  12.880 4.070 13.280 5.440 ;
        RECT  13.280 4.270 13.290 5.440 ;
        RECT  13.290 4.640 14.330 5.440 ;
        RECT  14.330 4.270 14.340 5.440 ;
        RECT  14.340 4.070 14.740 5.440 ;
        RECT  14.740 4.270 14.750 5.440 ;
        RECT  14.750 4.640 15.670 5.440 ;
        RECT  15.670 4.270 15.680 5.440 ;
        RECT  15.680 4.070 16.080 5.440 ;
        RECT  16.080 4.270 16.090 5.440 ;
        RECT  16.090 4.640 16.500 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        RECT  0.990 -0.400 1.390 0.560 ;
        RECT  1.390 -0.400 3.540 0.400 ;
        RECT  3.540 -0.400 3.940 1.310 ;
        RECT  3.940 -0.400 6.220 0.400 ;
        RECT  6.220 -0.400 6.230 1.200 ;
        RECT  6.230 -0.400 6.630 1.400 ;
        RECT  6.630 -0.400 6.640 1.200 ;
        RECT  6.640 -0.400 8.670 0.400 ;
        RECT  8.670 -0.400 9.070 1.310 ;
        RECT  9.070 -0.400 11.260 0.400 ;
        RECT  11.260 -0.400 11.660 0.560 ;
        RECT  11.660 -0.400 12.870 0.400 ;
        RECT  12.870 -0.400 12.880 0.730 ;
        RECT  12.880 -0.400 13.280 0.930 ;
        RECT  13.280 -0.400 13.290 0.730 ;
        RECT  13.290 -0.400 14.280 0.400 ;
        RECT  14.280 -0.400 14.290 1.010 ;
        RECT  14.290 -0.400 14.690 1.490 ;
        RECT  14.690 -0.400 14.700 1.010 ;
        RECT  14.700 -0.400 15.670 0.400 ;
        RECT  15.670 -0.400 15.680 0.730 ;
        RECT  15.680 -0.400 16.080 0.930 ;
        RECT  16.080 -0.400 16.090 0.730 ;
        RECT  16.090 -0.400 16.500 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  15.710 2.260 15.950 3.790 ;
        RECT  13.040 3.550 15.710 3.790 ;
        RECT  12.800 1.260 13.040 3.790 ;
        RECT  12.480 1.260 12.800 1.500 ;
        RECT  12.010 3.390 12.800 3.790 ;
        RECT  12.280 2.260 12.520 3.050 ;
        RECT  12.080 1.100 12.480 1.500 ;
        RECT  11.110 2.810 12.280 3.050 ;
        RECT  11.630 1.260 12.080 1.500 ;
        RECT  11.390 1.260 11.630 2.520 ;
        RECT  10.870 0.990 11.110 3.860 ;
        RECT  9.630 0.990 10.870 1.230 ;
        RECT  10.340 3.620 10.870 3.860 ;
        RECT  10.300 1.510 10.540 2.910 ;
        RECT  9.940 3.620 10.340 4.020 ;
        RECT  10.010 2.670 10.300 2.910 ;
        RECT  9.850 2.670 10.010 3.070 ;
        RECT  7.860 3.620 9.940 3.860 ;
        RECT  9.610 2.670 9.850 3.340 ;
        RECT  9.390 0.990 9.630 1.830 ;
        RECT  7.850 3.100 9.610 3.340 ;
        RECT  7.850 1.590 9.390 1.830 ;
        RECT  8.420 2.110 9.320 2.510 ;
        RECT  6.880 2.110 8.420 2.350 ;
        RECT  7.620 3.620 7.860 4.110 ;
        RECT  7.450 1.240 7.850 1.830 ;
        RECT  7.450 2.640 7.850 3.340 ;
        RECT  7.460 3.710 7.620 4.110 ;
        RECT  5.730 3.100 7.450 3.340 ;
        RECT  6.470 1.670 6.880 2.360 ;
        RECT  5.950 1.680 6.470 1.920 ;
        RECT  5.710 0.760 5.950 1.920 ;
        RECT  5.430 3.030 5.730 3.430 ;
        RECT  4.700 0.760 5.710 1.000 ;
        RECT  5.190 1.280 5.430 4.180 ;
        RECT  5.120 1.280 5.190 1.680 ;
        RECT  3.210 3.940 5.190 4.180 ;
        RECT  4.690 3.420 4.850 3.660 ;
        RECT  4.690 0.760 4.700 1.500 ;
        RECT  4.460 0.760 4.690 3.660 ;
        RECT  4.450 1.100 4.460 3.660 ;
        RECT  4.300 1.100 4.450 1.500 ;
        RECT  3.370 2.580 4.450 2.980 ;
        RECT  3.770 1.860 4.170 2.260 ;
        RECT  3.100 1.940 3.770 2.180 ;
        RECT  2.970 3.940 3.210 4.240 ;
        RECT  2.860 1.370 3.100 3.520 ;
        RECT  2.170 4.000 2.970 4.240 ;
        RECT  2.520 0.670 2.920 0.920 ;
        RECT  2.600 1.370 2.860 1.610 ;
        RECT  2.690 3.280 2.860 3.520 ;
        RECT  2.450 3.280 2.690 3.680 ;
        RECT  2.200 1.210 2.600 1.610 ;
        RECT  1.920 0.680 2.520 0.920 ;
        RECT  2.170 1.890 2.380 3.000 ;
        RECT  2.140 1.890 2.170 4.240 ;
        RECT  1.930 2.760 2.140 4.240 ;
        RECT  1.680 0.680 1.920 1.400 ;
        RECT  0.570 1.160 1.680 1.400 ;
        RECT  0.410 1.160 0.570 1.560 ;
        RECT  0.410 3.500 0.570 3.900 ;
        RECT  0.170 1.160 0.410 3.900 ;
    END
END DFFNX4

MACRO DFFNX2
    CLASS CORE ;
    FOREIGN DFFNX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.230 3.130 13.310 4.110 ;
        RECT  13.150 0.730 13.310 1.710 ;
        RECT  13.310 0.730 13.470 4.110 ;
        RECT  13.470 0.730 13.550 4.100 ;
        RECT  13.550 2.390 13.660 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.350 3.130 11.750 3.530 ;
        RECT  11.400 0.690 11.810 1.100 ;
        RECT  11.750 3.130 12.180 3.370 ;
        RECT  11.810 0.860 12.180 1.100 ;
        RECT  12.180 0.860 12.420 3.370 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.230 1.760 1.240 2.100 ;
        RECT  1.240 1.690 1.640 2.100 ;
        RECT  1.640 1.760 1.780 2.100 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.670 2.400 0.860 2.820 ;
        RECT  0.860 2.390 1.120 2.820 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 4.480 1.390 5.440 ;
        RECT  1.390 4.640 5.640 5.440 ;
        RECT  5.640 4.480 6.040 5.440 ;
        RECT  6.040 4.640 8.200 5.440 ;
        RECT  8.200 4.480 8.600 5.440 ;
        RECT  8.600 4.640 10.410 5.440 ;
        RECT  10.410 4.480 10.810 5.440 ;
        RECT  10.810 4.640 12.230 5.440 ;
        RECT  12.230 4.480 12.630 5.440 ;
        RECT  12.630 4.640 13.860 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        RECT  0.990 -0.400 1.390 0.560 ;
        RECT  1.390 -0.400 3.590 0.400 ;
        RECT  3.590 -0.400 3.600 1.220 ;
        RECT  3.600 -0.400 4.000 1.420 ;
        RECT  4.000 -0.400 4.010 1.220 ;
        RECT  4.010 -0.400 6.000 0.400 ;
        RECT  6.000 -0.400 6.400 1.400 ;
        RECT  6.400 -0.400 8.440 0.400 ;
        RECT  8.440 -0.400 8.840 1.400 ;
        RECT  8.840 -0.400 10.620 0.400 ;
        RECT  10.620 -0.400 10.630 0.790 ;
        RECT  10.630 -0.400 11.030 0.990 ;
        RECT  11.030 -0.400 11.040 0.790 ;
        RECT  11.040 -0.400 12.330 0.400 ;
        RECT  12.330 -0.400 12.730 0.560 ;
        RECT  12.730 -0.400 13.860 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.700 2.170 12.940 4.090 ;
        RECT  11.750 3.850 12.700 4.090 ;
        RECT  11.530 1.380 11.770 2.760 ;
        RECT  11.350 3.850 11.750 4.320 ;
        RECT  11.070 2.520 11.530 2.760 ;
        RECT  11.070 3.850 11.350 4.090 ;
        RECT  11.190 1.840 11.270 2.240 ;
        RECT  10.870 1.600 11.190 2.240 ;
        RECT  10.830 2.520 11.070 4.090 ;
        RECT  9.950 1.600 10.870 1.840 ;
        RECT  10.470 2.520 10.830 2.760 ;
        RECT  10.230 2.180 10.470 2.760 ;
        RECT  9.710 1.600 9.950 3.650 ;
        RECT  9.690 1.600 9.710 1.920 ;
        RECT  9.340 3.410 9.710 3.650 ;
        RECT  9.290 1.110 9.690 1.920 ;
        RECT  9.190 2.410 9.430 2.860 ;
        RECT  8.940 3.410 9.340 3.810 ;
        RECT  7.620 1.680 9.290 1.920 ;
        RECT  7.320 2.620 9.190 2.860 ;
        RECT  7.320 3.520 8.940 3.760 ;
        RECT  7.380 1.240 7.620 1.920 ;
        RECT  7.220 1.240 7.380 1.640 ;
        RECT  6.920 2.620 7.320 3.020 ;
        RECT  6.920 3.520 7.320 3.920 ;
        RECT  6.680 1.790 6.920 3.240 ;
        RECT  5.440 1.790 6.680 2.030 ;
        RECT  6.640 3.000 6.680 3.240 ;
        RECT  6.400 3.000 6.640 4.180 ;
        RECT  5.360 3.940 6.400 4.180 ;
        RECT  6.120 2.320 6.340 2.720 ;
        RECT  5.880 2.320 6.120 3.660 ;
        RECT  4.840 3.420 5.880 3.660 ;
        RECT  5.260 1.000 5.440 3.060 ;
        RECT  5.120 3.940 5.360 4.330 ;
        RECT  5.200 1.000 5.260 3.140 ;
        RECT  4.860 2.740 5.200 3.140 ;
        RECT  3.200 4.090 5.120 4.330 ;
        RECT  4.780 1.100 4.920 2.460 ;
        RECT  4.580 3.420 4.840 3.800 ;
        RECT  4.680 1.020 4.780 2.460 ;
        RECT  4.380 1.020 4.680 1.420 ;
        RECT  4.580 2.220 4.680 2.460 ;
        RECT  4.340 2.220 4.580 3.800 ;
        RECT  3.000 1.700 4.400 1.940 ;
        RECT  3.300 2.420 4.340 2.660 ;
        RECT  2.800 3.930 3.200 4.330 ;
        RECT  2.760 1.370 3.000 3.640 ;
        RECT  1.960 0.680 2.910 0.920 ;
        RECT  2.220 3.930 2.800 4.170 ;
        RECT  2.660 1.370 2.760 1.610 ;
        RECT  2.500 3.400 2.760 3.640 ;
        RECT  2.260 1.200 2.660 1.610 ;
        RECT  2.220 1.890 2.380 2.650 ;
        RECT  2.140 1.890 2.220 4.170 ;
        RECT  1.980 2.410 2.140 4.170 ;
        RECT  1.720 0.680 1.960 1.270 ;
        RECT  0.570 1.030 1.720 1.270 ;
        RECT  0.400 1.030 0.570 1.430 ;
        RECT  0.400 3.190 0.570 3.590 ;
        RECT  0.170 1.030 0.400 3.590 ;
        RECT  0.160 1.110 0.170 3.430 ;
    END
END DFFNX2

MACRO DFFNX1
    CLASS CORE ;
    FOREIGN DFFNX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFNXL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.310 1.320 11.330 1.720 ;
        RECT  11.330 1.320 11.710 3.410 ;
        RECT  11.710 1.430 11.720 3.410 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.760 3.130 10.160 3.530 ;
        RECT  9.870 0.690 10.440 1.100 ;
        RECT  10.160 3.130 10.790 3.370 ;
        RECT  10.440 0.860 10.790 1.100 ;
        RECT  10.790 0.860 11.030 3.370 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.670 1.890 2.320 ;
        END
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 0.870 2.650 ;
        RECT  0.870 2.390 1.120 3.030 ;
        RECT  1.120 2.630 1.510 3.030 ;
        END
    END CKN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.450 5.440 ;
        RECT  1.450 4.480 1.850 5.440 ;
        RECT  1.850 4.640 6.490 5.440 ;
        RECT  6.490 4.480 6.890 5.440 ;
        RECT  6.890 4.640 8.940 5.440 ;
        RECT  8.940 4.480 9.340 5.440 ;
        RECT  9.340 4.640 10.550 5.440 ;
        RECT  10.550 4.480 10.950 5.440 ;
        RECT  10.950 4.640 11.880 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.000 0.400 ;
        RECT  1.000 -0.400 1.410 0.410 ;
        RECT  1.410 -0.400 1.810 0.560 ;
        RECT  1.810 -0.400 4.100 0.400 ;
        RECT  4.100 -0.400 4.500 1.230 ;
        RECT  4.500 -0.400 6.650 0.400 ;
        RECT  6.650 -0.400 6.660 1.200 ;
        RECT  6.660 -0.400 7.060 1.400 ;
        RECT  7.060 -0.400 7.070 1.200 ;
        RECT  7.070 -0.400 9.100 0.400 ;
        RECT  9.100 -0.400 9.110 0.670 ;
        RECT  9.110 -0.400 9.510 0.870 ;
        RECT  9.510 -0.400 9.520 0.670 ;
        RECT  9.520 -0.400 10.720 0.400 ;
        RECT  10.720 -0.400 11.120 0.560 ;
        RECT  11.120 -0.400 11.880 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.310 1.430 10.550 2.830 ;
        RECT  9.930 1.430 10.310 1.670 ;
        RECT  9.070 2.590 10.310 2.830 ;
        RECT  9.760 3.940 10.160 4.360 ;
        RECT  9.610 2.000 9.800 2.240 ;
        RECT  9.050 3.940 9.760 4.180 ;
        RECT  9.370 1.600 9.610 2.240 ;
        RECT  8.380 1.600 9.370 1.840 ;
        RECT  9.050 2.130 9.070 2.830 ;
        RECT  8.810 2.130 9.050 4.180 ;
        RECT  8.670 2.130 8.810 2.530 ;
        RECT  7.600 0.760 8.610 1.000 ;
        RECT  8.280 1.440 8.380 3.940 ;
        RECT  8.170 1.280 8.280 3.940 ;
        RECT  8.140 1.280 8.170 4.100 ;
        RECT  7.880 1.280 8.140 1.680 ;
        RECT  7.770 3.700 8.140 4.100 ;
        RECT  7.600 2.480 7.830 2.880 ;
        RECT  7.490 0.760 7.600 2.880 ;
        RECT  7.360 0.760 7.490 4.180 ;
        RECT  7.250 1.800 7.360 4.180 ;
        RECT  6.180 1.800 7.250 2.040 ;
        RECT  6.210 3.940 7.250 4.180 ;
        RECT  6.730 2.320 6.970 3.660 ;
        RECT  5.690 3.420 6.730 3.660 ;
        RECT  5.970 3.940 6.210 4.370 ;
        RECT  6.020 1.280 6.180 2.040 ;
        RECT  5.780 1.280 6.020 3.140 ;
        RECT  4.120 4.130 5.970 4.370 ;
        RECT  5.620 2.740 5.780 3.140 ;
        RECT  5.450 3.420 5.690 3.850 ;
        RECT  4.860 3.610 5.450 3.850 ;
        RECT  5.220 0.980 5.380 1.380 ;
        RECT  4.980 0.980 5.220 2.390 ;
        RECT  4.860 2.150 4.980 2.390 ;
        RECT  4.600 2.150 4.860 3.850 ;
        RECT  3.870 1.510 4.700 1.750 ;
        RECT  4.220 2.150 4.600 2.550 ;
        RECT  3.880 2.830 4.120 4.370 ;
        RECT  2.920 2.830 3.880 3.070 ;
        RECT  3.500 3.910 3.880 4.370 ;
        RECT  3.630 1.500 3.870 1.750 ;
        RECT  3.160 1.500 3.630 1.740 ;
        RECT  2.400 3.340 3.580 3.580 ;
        RECT  2.780 3.910 3.180 4.310 ;
        RECT  2.760 1.070 3.160 1.740 ;
        RECT  2.680 2.020 2.920 3.070 ;
        RECT  1.030 3.910 2.780 4.150 ;
        RECT  2.400 1.500 2.760 1.740 ;
        RECT  2.160 1.500 2.400 3.580 ;
        RECT  0.790 3.320 1.030 4.150 ;
        RECT  0.530 1.110 0.930 1.510 ;
        RECT  0.630 3.320 0.790 3.720 ;
        RECT  0.500 3.320 0.630 3.560 ;
        RECT  0.500 1.270 0.530 1.510 ;
        RECT  0.260 1.270 0.500 3.560 ;
    END
END DFFNX1

MACRO DFFHQXL
    CLASS CORE ;
    FOREIGN DFFHQXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.380 3.250 9.440 3.510 ;
        RECT  9.440 3.250 9.700 3.770 ;
        RECT  9.700 3.250 9.790 3.510 ;
        RECT  9.790 3.250 10.160 3.490 ;
        RECT  9.560 0.640 10.160 0.880 ;
        RECT  10.160 0.640 10.400 3.490 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.390 1.760 2.930 ;
        RECT  1.760 2.390 1.780 2.920 ;
        RECT  1.780 2.400 1.990 2.920 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.760 2.940 0.770 3.290 ;
        RECT  0.770 2.860 1.010 3.290 ;
        RECT  1.010 2.940 1.210 3.290 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.520 5.440 ;
        RECT  1.520 4.390 1.530 5.440 ;
        RECT  1.530 4.270 1.930 5.440 ;
        RECT  1.930 4.390 1.940 5.440 ;
        RECT  1.940 4.640 4.150 5.440 ;
        RECT  4.150 4.390 4.160 5.440 ;
        RECT  4.160 4.270 4.560 5.440 ;
        RECT  4.560 4.390 4.570 5.440 ;
        RECT  4.570 4.640 6.450 5.440 ;
        RECT  6.450 4.480 6.850 5.440 ;
        RECT  6.850 4.640 8.130 5.440 ;
        RECT  8.130 4.480 8.530 5.440 ;
        RECT  8.530 4.640 10.560 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.040 0.400 ;
        RECT  1.040 -0.400 1.440 0.560 ;
        RECT  1.440 -0.400 3.300 0.400 ;
        RECT  3.300 -0.400 3.310 0.730 ;
        RECT  3.310 -0.400 3.710 0.930 ;
        RECT  3.710 -0.400 3.720 0.730 ;
        RECT  3.720 -0.400 5.660 0.400 ;
        RECT  5.660 -0.400 5.670 0.730 ;
        RECT  5.670 -0.400 6.070 0.930 ;
        RECT  6.070 -0.400 6.080 0.730 ;
        RECT  6.080 -0.400 8.640 0.400 ;
        RECT  8.640 -0.400 8.650 0.670 ;
        RECT  8.650 -0.400 9.050 0.870 ;
        RECT  9.050 -0.400 9.060 0.670 ;
        RECT  9.060 -0.400 10.560 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  9.640 1.330 9.880 2.970 ;
        RECT  9.050 4.030 9.780 4.270 ;
        RECT  8.630 2.730 9.640 2.970 ;
        RECT  9.120 1.350 9.360 2.450 ;
        RECT  8.110 1.350 9.120 1.590 ;
        RECT  8.810 3.940 9.050 4.270 ;
        RECT  8.630 3.940 8.810 4.180 ;
        RECT  8.390 2.110 8.630 4.180 ;
        RECT  7.360 0.680 8.280 0.920 ;
        RECT  7.880 1.350 8.110 3.750 ;
        RECT  7.870 1.200 7.880 3.750 ;
        RECT  7.640 1.200 7.870 1.600 ;
        RECT  7.360 2.000 7.590 4.260 ;
        RECT  7.350 0.680 7.360 4.260 ;
        RECT  7.120 0.680 7.350 2.240 ;
        RECT  7.150 3.940 7.350 4.260 ;
        RECT  6.150 3.940 7.150 4.180 ;
        RECT  6.840 2.520 7.060 3.200 ;
        RECT  6.820 1.330 6.840 3.200 ;
        RECT  6.810 1.330 6.820 2.760 ;
        RECT  6.600 1.170 6.810 2.760 ;
        RECT  6.570 1.170 6.600 1.570 ;
        RECT  6.080 1.850 6.320 3.470 ;
        RECT  5.910 3.940 6.150 4.370 ;
        RECT  5.600 3.230 6.080 3.470 ;
        RECT  5.080 4.130 5.910 4.370 ;
        RECT  5.360 3.230 5.600 3.840 ;
        RECT  5.170 2.680 5.380 2.920 ;
        RECT  4.590 3.230 5.360 3.470 ;
        RECT  5.170 1.170 5.330 1.570 ;
        RECT  4.930 0.670 5.170 2.920 ;
        RECT  4.840 3.750 5.080 4.370 ;
        RECT  4.330 0.670 4.930 0.910 ;
        RECT  3.810 3.750 4.840 3.990 ;
        RECT  4.350 1.250 4.590 3.470 ;
        RECT  4.190 1.250 4.350 1.490 ;
        RECT  4.220 2.630 4.350 3.470 ;
        RECT  3.930 2.630 4.220 2.870 ;
        RECT  3.390 1.830 4.070 2.070 ;
        RECT  3.690 2.470 3.930 2.870 ;
        RECT  3.370 3.750 3.810 4.350 ;
        RECT  3.150 1.830 3.390 3.470 ;
        RECT  2.510 3.750 3.370 3.990 ;
        RECT  3.030 1.830 3.150 2.070 ;
        RECT  2.790 1.160 3.030 2.070 ;
        RECT  2.190 1.160 2.790 1.400 ;
        RECT  2.270 1.830 2.510 3.990 ;
        RECT  2.050 1.830 2.270 2.070 ;
        RECT  0.480 3.560 2.270 3.800 ;
        RECT  0.480 1.060 0.570 1.460 ;
        RECT  0.240 1.060 0.480 3.800 ;
        RECT  0.170 1.060 0.240 1.460 ;
    END
END DFFHQXL

MACRO DFFHQX4
    CLASS CORE ;
    FOREIGN DFFHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFHQXL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.690 0.660 13.850 1.640 ;
        RECT  13.710 2.730 13.970 3.740 ;
        RECT  13.850 0.660 13.970 2.060 ;
        RECT  13.970 0.660 14.090 3.740 ;
        RECT  14.090 1.820 14.110 3.740 ;
        RECT  14.110 1.820 14.410 3.220 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.250 1.260 1.870 1.590 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.720 1.970 0.860 2.640 ;
        RECT  0.860 1.970 0.960 2.650 ;
        RECT  0.960 2.390 1.120 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.070 5.440 ;
        RECT  1.070 4.480 1.470 5.440 ;
        RECT  1.470 4.640 3.530 5.440 ;
        RECT  3.530 4.480 3.930 5.440 ;
        RECT  3.930 4.640 5.870 5.440 ;
        RECT  5.870 4.050 5.880 5.440 ;
        RECT  5.880 3.930 6.280 5.440 ;
        RECT  6.280 4.050 6.290 5.440 ;
        RECT  6.290 4.640 9.640 5.440 ;
        RECT  9.640 3.980 9.650 5.440 ;
        RECT  9.650 3.860 10.050 5.440 ;
        RECT  10.050 3.980 10.060 5.440 ;
        RECT  10.060 4.640 11.420 5.440 ;
        RECT  11.420 4.480 11.820 5.440 ;
        RECT  11.820 4.640 13.130 5.440 ;
        RECT  12.950 3.300 13.130 3.700 ;
        RECT  13.130 3.300 13.370 5.440 ;
        RECT  13.370 4.640 14.530 5.440 ;
        RECT  14.530 3.820 14.930 5.440 ;
        RECT  14.930 4.640 15.180 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.000 0.400 ;
        RECT  1.000 -0.400 1.400 0.970 ;
        RECT  1.400 -0.400 3.390 0.400 ;
        RECT  3.390 -0.400 3.400 0.750 ;
        RECT  3.400 -0.400 3.800 0.870 ;
        RECT  3.800 -0.400 3.810 0.750 ;
        RECT  3.810 -0.400 5.890 0.400 ;
        RECT  5.890 -0.400 5.900 1.080 ;
        RECT  5.900 -0.400 6.300 1.200 ;
        RECT  6.300 -0.400 6.310 1.080 ;
        RECT  6.310 -0.400 9.750 0.400 ;
        RECT  9.750 -0.400 10.150 0.560 ;
        RECT  10.150 -0.400 11.300 0.400 ;
        RECT  11.300 -0.400 11.700 0.560 ;
        RECT  11.700 -0.400 12.920 0.400 ;
        RECT  12.920 -0.400 12.930 0.980 ;
        RECT  12.930 -0.400 13.330 1.470 ;
        RECT  13.330 -0.400 13.340 0.980 ;
        RECT  13.340 -0.400 14.500 0.400 ;
        RECT  14.500 -0.400 14.510 1.020 ;
        RECT  14.510 -0.400 14.910 1.220 ;
        RECT  14.910 -0.400 14.920 1.020 ;
        RECT  14.920 -0.400 14.930 0.560 ;
        RECT  14.930 -0.400 15.180 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.650 4.130 12.850 4.370 ;
        RECT  12.410 1.150 12.650 4.370 ;
        RECT  12.170 1.150 12.410 1.390 ;
        RECT  11.690 2.470 12.410 2.870 ;
        RECT  11.910 1.630 12.130 2.030 ;
        RECT  11.490 1.630 11.910 2.040 ;
        RECT  11.450 1.190 11.490 2.040 ;
        RECT  11.210 1.190 11.450 3.070 ;
        RECT  10.570 1.190 11.210 1.430 ;
        RECT  10.920 2.830 11.210 3.070 ;
        RECT  10.730 1.710 10.970 2.550 ;
        RECT  8.900 1.710 10.730 1.950 ;
        RECT  10.170 1.140 10.570 1.430 ;
        RECT  8.220 1.190 10.170 1.430 ;
        RECT  9.500 2.260 9.760 2.500 ;
        RECT  9.370 2.260 9.500 3.580 ;
        RECT  9.260 2.260 9.370 4.120 ;
        RECT  7.700 0.670 9.290 0.910 ;
        RECT  9.130 3.340 9.260 4.120 ;
        RECT  6.800 3.880 9.130 4.120 ;
        RECT  8.840 2.660 8.980 3.060 ;
        RECT  8.500 1.710 8.900 2.030 ;
        RECT  8.600 2.660 8.840 3.600 ;
        RECT  7.700 3.360 8.600 3.600 ;
        RECT  7.980 1.190 8.220 3.080 ;
        RECT  7.460 0.670 7.700 3.600 ;
        RECT  6.660 0.670 7.460 0.910 ;
        RECT  7.140 2.690 7.460 3.090 ;
        RECT  6.940 1.480 7.180 2.130 ;
        RECT  5.410 1.480 6.940 1.720 ;
        RECT  6.560 3.190 6.800 4.120 ;
        RECT  6.360 3.190 6.560 3.430 ;
        RECT  6.120 2.000 6.360 3.430 ;
        RECT  4.730 3.190 6.120 3.430 ;
        RECT  3.240 3.710 5.600 3.950 ;
        RECT  5.250 2.650 5.480 2.890 ;
        RECT  5.250 1.190 5.410 1.720 ;
        RECT  5.010 0.680 5.250 2.890 ;
        RECT  4.550 0.680 5.010 0.920 ;
        RECT  4.490 1.270 4.730 3.430 ;
        RECT  4.220 1.270 4.490 1.510 ;
        RECT  3.510 3.190 4.490 3.430 ;
        RECT  3.790 1.840 4.190 2.100 ;
        RECT  2.720 1.840 3.790 2.080 ;
        RECT  3.270 2.400 3.510 3.430 ;
        RECT  3.040 2.400 3.270 2.640 ;
        RECT  3.000 3.710 3.240 4.160 ;
        RECT  2.120 3.920 3.000 4.160 ;
        RECT  2.480 1.040 2.720 3.610 ;
        RECT  2.360 1.040 2.480 1.440 ;
        RECT  1.880 2.060 2.120 4.160 ;
        RECT  0.640 3.310 1.880 3.550 ;
        RECT  0.410 3.300 0.640 4.320 ;
        RECT  0.410 0.930 0.570 1.330 ;
        RECT  0.240 0.930 0.410 4.320 ;
        RECT  0.170 0.930 0.240 3.540 ;
    END
END DFFHQX4

MACRO DFFHQX2
    CLASS CORE ;
    FOREIGN DFFHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFHQXL ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.000 2.920 11.240 3.320 ;
        RECT  11.240 2.920 11.340 3.220 ;
        RECT  11.340 1.280 11.420 3.220 ;
        RECT  11.420 1.270 11.430 3.220 ;
        RECT  11.430 1.270 11.580 3.160 ;
        RECT  11.580 1.270 11.680 1.530 ;
        RECT  11.680 1.270 11.740 1.510 ;
        RECT  11.740 0.930 12.140 1.510 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 1.820 1.630 2.100 ;
        RECT  1.630 1.820 1.870 2.350 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.770 2.380 1.220 2.800 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.720 5.440 ;
        RECT  1.720 3.920 1.730 5.440 ;
        RECT  1.730 3.800 2.130 5.440 ;
        RECT  2.130 3.920 2.140 5.440 ;
        RECT  2.140 4.640 4.040 5.440 ;
        RECT  4.040 4.390 4.050 5.440 ;
        RECT  4.050 4.270 4.450 5.440 ;
        RECT  4.450 4.390 4.460 5.440 ;
        RECT  4.460 4.640 6.110 5.440 ;
        RECT  6.110 4.160 6.510 5.440 ;
        RECT  6.510 4.640 9.960 5.440 ;
        RECT  9.960 3.240 10.200 5.440 ;
        RECT  10.200 4.640 11.730 5.440 ;
        RECT  11.730 3.790 11.740 5.440 ;
        RECT  11.740 3.590 12.140 5.440 ;
        RECT  12.140 3.790 12.150 5.440 ;
        RECT  12.150 4.640 12.540 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.300 0.400 ;
        RECT  0.300 -0.400 0.700 0.560 ;
        RECT  0.700 -0.400 3.300 0.400 ;
        RECT  3.300 -0.400 3.310 0.730 ;
        RECT  3.310 -0.400 3.710 0.930 ;
        RECT  3.710 -0.400 3.720 0.730 ;
        RECT  3.720 -0.400 5.810 0.400 ;
        RECT  5.810 -0.400 6.210 0.560 ;
        RECT  6.210 -0.400 9.600 0.400 ;
        RECT  9.600 -0.400 10.000 0.560 ;
        RECT  10.000 -0.400 10.910 0.400 ;
        RECT  10.910 -0.400 11.310 0.560 ;
        RECT  11.310 -0.400 12.540 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.760 3.850 11.160 4.250 ;
        RECT  10.720 1.130 10.790 2.640 ;
        RECT  10.720 3.850 10.760 4.090 ;
        RECT  10.550 1.130 10.720 4.090 ;
        RECT  10.480 2.400 10.550 4.090 ;
        RECT  9.400 2.400 10.480 2.640 ;
        RECT  10.030 1.230 10.270 2.120 ;
        RECT  8.790 1.230 10.030 1.470 ;
        RECT  7.030 4.110 9.680 4.350 ;
        RECT  9.160 2.090 9.400 2.640 ;
        RECT  9.070 3.300 9.310 3.830 ;
        RECT  6.730 0.670 9.170 0.910 ;
        RECT  7.550 3.590 9.070 3.830 ;
        RECT  8.550 1.190 8.790 3.280 ;
        RECT  7.990 3.040 8.550 3.280 ;
        RECT  8.030 1.190 8.270 2.700 ;
        RECT  7.010 1.190 8.030 1.430 ;
        RECT  7.550 2.460 8.030 2.700 ;
        RECT  7.510 1.710 7.750 2.160 ;
        RECT  7.310 2.460 7.550 3.830 ;
        RECT  6.470 1.710 7.510 1.950 ;
        RECT  6.790 2.320 7.030 4.350 ;
        RECT  5.490 3.610 6.790 3.850 ;
        RECT  6.490 0.670 6.730 1.110 ;
        RECT  5.950 0.870 6.490 1.110 ;
        RECT  6.230 1.710 6.470 2.920 ;
        RECT  6.010 2.680 6.230 2.920 ;
        RECT  5.770 2.680 6.010 3.080 ;
        RECT  5.710 0.870 5.950 2.290 ;
        RECT  4.970 4.130 5.800 4.370 ;
        RECT  5.110 2.680 5.770 2.920 ;
        RECT  5.250 3.230 5.490 3.850 ;
        RECT  5.110 1.170 5.430 1.590 ;
        RECT  4.590 3.230 5.250 3.470 ;
        RECT  4.870 0.670 5.110 2.920 ;
        RECT  4.730 3.750 4.970 4.370 ;
        RECT  4.300 0.670 4.870 0.910 ;
        RECT  3.770 3.750 4.730 3.990 ;
        RECT  4.350 1.260 4.590 3.470 ;
        RECT  4.190 1.260 4.350 1.500 ;
        RECT  3.900 2.460 4.350 2.870 ;
        RECT  3.390 1.830 4.070 2.070 ;
        RECT  3.690 2.470 3.900 2.870 ;
        RECT  3.530 3.750 3.770 4.350 ;
        RECT  2.670 4.110 3.530 4.350 ;
        RECT  3.150 1.830 3.390 3.470 ;
        RECT  2.910 1.830 3.150 2.070 ;
        RECT  2.670 0.750 2.910 2.070 ;
        RECT  2.190 0.750 2.670 0.990 ;
        RECT  2.430 3.280 2.670 4.350 ;
        RECT  2.390 3.280 2.430 3.520 ;
        RECT  2.150 1.310 2.390 3.520 ;
        RECT  1.810 1.310 2.150 1.550 ;
        RECT  1.220 3.280 2.150 3.520 ;
        RECT  0.820 3.280 1.220 3.680 ;
        RECT  0.500 3.280 0.820 3.520 ;
        RECT  0.500 1.290 0.570 1.690 ;
        RECT  0.260 1.290 0.500 3.520 ;
        RECT  0.170 1.290 0.260 1.690 ;
    END
END DFFHQX2

MACRO DFFHQX1
    CLASS CORE ;
    FOREIGN DFFHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFHQXL ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.320 3.250 9.350 3.490 ;
        RECT  9.350 3.250 9.440 3.510 ;
        RECT  9.440 3.250 9.700 3.770 ;
        RECT  9.700 3.250 9.790 3.510 ;
        RECT  9.790 3.250 10.160 3.490 ;
        RECT  9.500 0.670 10.160 0.910 ;
        RECT  10.160 0.670 10.400 3.490 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.330 1.880 1.530 2.280 ;
        RECT  1.520 1.270 1.530 1.530 ;
        RECT  1.530 1.270 1.770 2.280 ;
        RECT  1.770 1.270 1.780 1.530 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.770 2.750 1.320 3.220 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.540 5.440 ;
        RECT  1.540 4.390 1.550 5.440 ;
        RECT  1.550 4.270 1.950 5.440 ;
        RECT  1.950 4.390 1.960 5.440 ;
        RECT  1.960 4.640 4.150 5.440 ;
        RECT  4.150 4.390 4.160 5.440 ;
        RECT  4.160 4.270 4.560 5.440 ;
        RECT  4.560 4.390 4.570 5.440 ;
        RECT  4.570 4.640 6.450 5.440 ;
        RECT  6.450 4.480 6.850 5.440 ;
        RECT  6.850 4.640 8.130 5.440 ;
        RECT  8.130 4.480 8.530 5.440 ;
        RECT  8.530 4.640 10.560 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.220 0.400 ;
        RECT  1.220 -0.400 1.620 0.560 ;
        RECT  1.620 -0.400 3.300 0.400 ;
        RECT  3.300 -0.400 3.310 0.730 ;
        RECT  3.310 -0.400 3.710 0.930 ;
        RECT  3.710 -0.400 3.720 0.730 ;
        RECT  3.720 -0.400 5.660 0.400 ;
        RECT  5.660 -0.400 5.670 0.730 ;
        RECT  5.670 -0.400 6.070 0.930 ;
        RECT  6.070 -0.400 6.080 0.730 ;
        RECT  6.080 -0.400 8.640 0.400 ;
        RECT  8.640 -0.400 8.650 0.670 ;
        RECT  8.650 -0.400 9.050 0.870 ;
        RECT  9.050 -0.400 9.060 0.670 ;
        RECT  9.060 -0.400 10.560 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  9.640 1.350 9.880 2.970 ;
        RECT  9.050 4.030 9.780 4.270 ;
        RECT  8.630 2.730 9.640 2.970 ;
        RECT  9.120 1.350 9.360 2.450 ;
        RECT  8.110 1.350 9.120 1.590 ;
        RECT  8.810 3.940 9.050 4.270 ;
        RECT  8.630 3.940 8.810 4.180 ;
        RECT  8.390 2.080 8.630 4.180 ;
        RECT  7.360 0.680 8.280 0.920 ;
        RECT  7.880 1.350 8.110 3.760 ;
        RECT  7.870 1.200 7.880 3.760 ;
        RECT  7.640 1.200 7.870 1.600 ;
        RECT  7.360 2.000 7.590 4.260 ;
        RECT  7.350 0.680 7.360 4.260 ;
        RECT  7.120 0.680 7.350 2.240 ;
        RECT  7.150 3.940 7.350 4.260 ;
        RECT  6.150 3.940 7.150 4.180 ;
        RECT  6.840 2.520 7.060 3.430 ;
        RECT  6.820 1.050 6.840 3.430 ;
        RECT  6.600 1.050 6.820 2.760 ;
        RECT  6.570 1.050 6.600 1.450 ;
        RECT  6.080 2.070 6.320 3.470 ;
        RECT  5.910 3.940 6.150 4.370 ;
        RECT  5.600 3.230 6.080 3.470 ;
        RECT  5.080 4.130 5.910 4.370 ;
        RECT  5.360 3.230 5.600 3.840 ;
        RECT  5.170 2.680 5.380 2.920 ;
        RECT  4.590 3.230 5.360 3.470 ;
        RECT  5.170 1.210 5.330 1.610 ;
        RECT  4.930 0.670 5.170 2.920 ;
        RECT  4.840 3.750 5.080 4.370 ;
        RECT  4.330 0.670 4.930 0.910 ;
        RECT  3.770 3.750 4.840 3.990 ;
        RECT  4.350 1.250 4.590 3.470 ;
        RECT  4.190 1.250 4.350 1.490 ;
        RECT  4.220 2.630 4.350 3.470 ;
        RECT  3.930 2.630 4.220 2.870 ;
        RECT  3.390 1.830 4.070 2.070 ;
        RECT  3.690 2.470 3.930 2.870 ;
        RECT  3.370 3.750 3.770 4.350 ;
        RECT  3.150 1.830 3.390 3.470 ;
        RECT  2.870 3.750 3.370 3.990 ;
        RECT  3.030 1.830 3.150 2.070 ;
        RECT  2.790 0.740 3.030 2.070 ;
        RECT  2.380 3.550 2.870 3.990 ;
        RECT  2.190 0.740 2.790 0.980 ;
        RECT  2.370 2.460 2.380 3.990 ;
        RECT  2.140 1.880 2.370 3.990 ;
        RECT  2.130 1.880 2.140 2.700 ;
        RECT  0.500 3.550 2.140 3.790 ;
        RECT  0.500 1.310 0.680 1.710 ;
        RECT  0.260 1.310 0.500 3.790 ;
    END
END DFFHQX1

MACRO DFFXL
    CLASS CORE ;
    FOREIGN DFFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.330 1.780 11.340 3.250 ;
        RECT  11.340 1.390 11.670 3.250 ;
        RECT  11.670 1.780 11.680 3.250 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.750 2.920 10.150 3.320 ;
        RECT  10.150 2.930 10.360 3.210 ;
        RECT  10.140 0.720 10.540 1.100 ;
        RECT  10.360 2.930 10.820 3.170 ;
        RECT  10.540 0.860 10.820 1.100 ;
        RECT  10.820 0.860 11.060 3.170 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.520 1.900 2.090 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.360 1.630 2.780 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.730 5.440 ;
        RECT  1.730 4.480 2.130 5.440 ;
        RECT  2.130 4.640 6.490 5.440 ;
        RECT  6.490 4.480 6.890 5.440 ;
        RECT  6.890 4.640 8.930 5.440 ;
        RECT  8.930 4.480 9.330 5.440 ;
        RECT  9.330 4.640 10.550 5.440 ;
        RECT  10.550 4.480 10.950 5.440 ;
        RECT  10.950 4.640 11.880 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.380 0.400 ;
        RECT  1.380 -0.400 1.780 0.560 ;
        RECT  1.780 -0.400 4.070 0.400 ;
        RECT  4.070 -0.400 4.470 1.180 ;
        RECT  4.470 -0.400 6.650 0.400 ;
        RECT  6.650 -0.400 6.660 1.380 ;
        RECT  6.660 -0.400 7.060 1.500 ;
        RECT  7.060 -0.400 7.070 1.380 ;
        RECT  7.070 -0.400 9.250 0.400 ;
        RECT  9.250 -0.400 9.260 0.880 ;
        RECT  9.260 -0.400 9.660 1.080 ;
        RECT  9.660 -0.400 9.670 0.880 ;
        RECT  9.670 -0.400 11.090 0.400 ;
        RECT  11.090 -0.400 11.490 0.560 ;
        RECT  11.490 -0.400 11.880 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.300 1.460 10.540 2.640 ;
        RECT  10.140 1.460 10.300 1.700 ;
        RECT  9.100 2.400 10.300 2.640 ;
        RECT  9.810 3.800 10.210 4.200 ;
        RECT  9.700 1.860 9.860 2.100 ;
        RECT  9.060 3.800 9.810 4.040 ;
        RECT  9.460 1.610 9.700 2.100 ;
        RECT  8.380 1.610 9.460 1.850 ;
        RECT  9.060 2.310 9.100 2.710 ;
        RECT  8.820 2.310 9.060 4.040 ;
        RECT  8.700 2.310 8.820 2.710 ;
        RECT  7.600 0.760 8.610 1.000 ;
        RECT  8.140 1.290 8.380 4.220 ;
        RECT  7.880 1.290 8.140 1.690 ;
        RECT  7.830 3.820 8.140 4.220 ;
        RECT  7.600 2.610 7.830 3.010 ;
        RECT  7.550 0.760 7.600 3.010 ;
        RECT  7.360 0.760 7.550 4.180 ;
        RECT  6.310 1.800 7.360 2.040 ;
        RECT  7.310 2.770 7.360 4.180 ;
        RECT  6.210 3.940 7.310 4.180 ;
        RECT  6.790 2.320 7.030 3.660 ;
        RECT  5.690 3.420 6.790 3.660 ;
        RECT  6.070 1.800 6.310 2.460 ;
        RECT  5.970 3.940 6.210 4.370 ;
        RECT  6.040 1.260 6.180 1.500 ;
        RECT  5.790 2.740 6.090 3.140 ;
        RECT  5.790 0.670 6.040 1.500 ;
        RECT  4.120 4.130 5.970 4.370 ;
        RECT  5.690 0.670 5.790 3.140 ;
        RECT  5.550 0.670 5.690 3.060 ;
        RECT  5.450 3.420 5.690 3.850 ;
        RECT  4.860 3.610 5.450 3.850 ;
        RECT  5.030 1.010 5.270 2.390 ;
        RECT  4.860 2.150 5.030 2.390 ;
        RECT  4.600 2.150 4.860 3.850 ;
        RECT  3.840 1.510 4.750 1.750 ;
        RECT  4.220 2.150 4.600 2.550 ;
        RECT  3.940 2.890 4.120 4.370 ;
        RECT  3.880 2.350 3.940 4.370 ;
        RECT  3.700 2.350 3.880 3.130 ;
        RECT  3.480 3.930 3.880 4.370 ;
        RECT  3.600 1.500 3.840 1.750 ;
        RECT  2.930 2.350 3.700 2.590 ;
        RECT  3.130 1.500 3.600 1.740 ;
        RECT  2.410 3.410 3.560 3.650 ;
        RECT  1.250 3.930 3.480 4.170 ;
        RECT  2.730 0.960 3.130 1.740 ;
        RECT  2.690 2.020 2.930 2.590 ;
        RECT  2.410 1.500 2.730 1.740 ;
        RECT  2.170 1.500 2.410 3.650 ;
        RECT  1.010 3.130 1.250 4.170 ;
        RECT  0.850 3.130 1.010 3.530 ;
        RECT  0.530 1.120 0.900 1.520 ;
        RECT  0.530 3.130 0.850 3.370 ;
        RECT  0.290 1.120 0.530 3.370 ;
    END
END DFFXL

MACRO DFFX4
    CLASS CORE ;
    FOREIGN DFFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  15.290 1.820 15.680 3.220 ;
        RECT  15.680 1.410 15.690 3.220 ;
        RECT  15.690 1.210 16.090 3.270 ;
        RECT  16.090 1.410 16.100 3.070 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.970 1.820 14.140 3.220 ;
        RECT  14.140 1.410 14.150 3.220 ;
        RECT  14.150 1.210 14.550 3.270 ;
        RECT  14.550 1.410 14.560 3.070 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.500 1.650 1.870 2.240 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.830 2.080 1.170 2.740 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.510 5.440 ;
        RECT  1.510 4.480 1.910 5.440 ;
        RECT  1.910 4.640 4.290 5.440 ;
        RECT  4.290 4.480 4.690 5.440 ;
        RECT  4.690 4.640 6.840 5.440 ;
        RECT  6.840 4.480 7.240 5.440 ;
        RECT  7.240 4.640 9.340 5.440 ;
        RECT  9.340 4.140 9.740 5.440 ;
        RECT  9.740 4.640 11.920 5.440 ;
        RECT  11.920 4.480 12.320 5.440 ;
        RECT  12.320 4.640 13.480 5.440 ;
        RECT  13.480 4.270 13.490 5.440 ;
        RECT  13.490 4.070 13.890 5.440 ;
        RECT  13.890 4.270 13.900 5.440 ;
        RECT  13.900 4.640 14.970 5.440 ;
        RECT  14.970 4.270 14.980 5.440 ;
        RECT  14.980 4.070 15.380 5.440 ;
        RECT  15.380 4.270 15.390 5.440 ;
        RECT  15.390 4.640 16.350 5.440 ;
        RECT  16.350 4.270 16.360 5.440 ;
        RECT  16.360 4.070 16.760 5.440 ;
        RECT  16.760 4.270 16.770 5.440 ;
        RECT  16.770 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.330 0.400 ;
        RECT  1.330 -0.400 1.340 0.890 ;
        RECT  1.340 -0.400 1.740 1.090 ;
        RECT  1.740 -0.400 1.750 0.890 ;
        RECT  1.750 -0.400 4.040 0.400 ;
        RECT  4.040 -0.400 4.440 1.300 ;
        RECT  4.440 -0.400 6.880 0.400 ;
        RECT  6.880 -0.400 6.890 1.200 ;
        RECT  6.890 -0.400 7.290 1.400 ;
        RECT  7.290 -0.400 7.300 1.200 ;
        RECT  7.300 -0.400 9.330 0.400 ;
        RECT  9.330 -0.400 9.730 1.300 ;
        RECT  9.730 -0.400 11.920 0.400 ;
        RECT  11.920 -0.400 12.320 0.560 ;
        RECT  12.320 -0.400 13.550 0.400 ;
        RECT  13.550 -0.400 13.560 0.730 ;
        RECT  13.560 -0.400 13.960 0.930 ;
        RECT  13.960 -0.400 13.970 0.730 ;
        RECT  13.970 -0.400 14.940 0.400 ;
        RECT  14.940 -0.400 14.950 1.010 ;
        RECT  14.950 -0.400 15.350 1.490 ;
        RECT  15.350 -0.400 15.360 1.010 ;
        RECT  15.360 -0.400 16.350 0.400 ;
        RECT  16.350 -0.400 16.360 0.730 ;
        RECT  16.360 -0.400 16.760 0.930 ;
        RECT  16.760 -0.400 16.770 0.730 ;
        RECT  16.770 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.430 2.260 16.670 3.790 ;
        RECT  13.700 3.550 16.430 3.790 ;
        RECT  13.460 1.260 13.700 3.790 ;
        RECT  13.140 1.260 13.460 1.500 ;
        RECT  12.690 3.390 13.460 3.790 ;
        RECT  12.940 2.260 13.180 3.050 ;
        RECT  12.740 1.100 13.140 1.500 ;
        RECT  11.770 2.810 12.940 3.050 ;
        RECT  12.290 1.260 12.740 1.500 ;
        RECT  12.050 1.260 12.290 2.520 ;
        RECT  11.530 1.000 11.770 3.860 ;
        RECT  10.290 1.000 11.530 1.240 ;
        RECT  11.000 3.620 11.530 3.860 ;
        RECT  10.960 1.510 11.200 2.910 ;
        RECT  10.600 3.620 11.000 4.020 ;
        RECT  10.760 2.670 10.960 2.910 ;
        RECT  10.360 2.670 10.760 3.340 ;
        RECT  8.520 3.620 10.600 3.860 ;
        RECT  8.320 3.100 10.360 3.340 ;
        RECT  10.050 1.000 10.290 1.830 ;
        RECT  8.510 1.590 10.050 1.830 ;
        RECT  9.090 2.110 9.490 2.510 ;
        RECT  7.540 2.110 9.090 2.350 ;
        RECT  8.200 3.620 8.520 4.110 ;
        RECT  8.110 1.240 8.510 1.830 ;
        RECT  7.920 2.640 8.320 3.340 ;
        RECT  8.120 3.710 8.200 4.110 ;
        RECT  7.840 3.100 7.920 3.340 ;
        RECT  7.600 3.100 7.840 4.180 ;
        RECT  6.830 3.940 7.600 4.180 ;
        RECT  7.460 1.920 7.540 2.630 ;
        RECT  7.130 1.680 7.460 2.630 ;
        RECT  6.610 1.680 7.130 1.920 ;
        RECT  6.590 2.210 6.830 4.180 ;
        RECT  6.370 0.760 6.610 1.920 ;
        RECT  6.400 2.210 6.590 2.610 ;
        RECT  3.870 3.940 6.590 4.180 ;
        RECT  5.200 0.760 6.370 1.000 ;
        RECT  6.090 3.030 6.310 3.430 ;
        RECT  5.850 1.280 6.090 3.430 ;
        RECT  5.690 1.280 5.850 2.260 ;
        RECT  5.490 1.860 5.690 2.260 ;
        RECT  5.200 3.420 5.510 3.660 ;
        RECT  4.960 0.760 5.200 3.660 ;
        RECT  4.800 1.100 4.960 1.500 ;
        RECT  4.550 2.660 4.960 2.900 ;
        RECT  4.280 1.830 4.680 2.180 ;
        RECT  4.150 2.580 4.550 2.980 ;
        RECT  3.430 1.830 4.280 2.070 ;
        RECT  3.630 2.350 3.870 4.240 ;
        RECT  2.900 2.350 3.630 2.590 ;
        RECT  2.600 4.000 3.630 4.240 ;
        RECT  3.190 1.420 3.430 2.070 ;
        RECT  3.110 3.310 3.350 3.710 ;
        RECT  3.070 1.420 3.190 1.660 ;
        RECT  2.380 3.310 3.110 3.550 ;
        RECT  2.670 0.690 3.070 1.660 ;
        RECT  2.660 1.940 2.900 2.590 ;
        RECT  2.380 1.420 2.670 1.660 ;
        RECT  2.360 3.840 2.600 4.240 ;
        RECT  2.140 1.420 2.380 3.550 ;
        RECT  1.090 3.840 2.360 4.080 ;
        RECT  0.690 3.110 1.090 4.090 ;
        RECT  0.520 0.890 0.920 1.290 ;
        RECT  0.500 3.110 0.690 3.350 ;
        RECT  0.500 1.050 0.520 1.290 ;
        RECT  0.260 1.050 0.500 3.350 ;
    END
END DFFX4

MACRO DFFX2
    CLASS CORE ;
    FOREIGN DFFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFXL ;
    SIZE 14.520 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.890 3.130 13.970 4.110 ;
        RECT  13.810 0.730 13.970 1.710 ;
        RECT  13.970 0.730 14.130 4.110 ;
        RECT  14.130 0.730 14.210 4.100 ;
        RECT  14.210 2.390 14.320 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.060 0.690 12.470 1.100 ;
        RECT  12.010 3.130 12.840 3.530 ;
        RECT  12.470 0.860 12.840 1.100 ;
        RECT  12.840 0.860 13.080 3.530 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.700 1.870 2.230 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.840 1.980 1.150 2.650 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.670 5.440 ;
        RECT  1.670 4.480 2.070 5.440 ;
        RECT  2.070 4.640 6.300 5.440 ;
        RECT  6.300 4.480 6.700 5.440 ;
        RECT  6.700 4.640 8.860 5.440 ;
        RECT  8.860 4.480 9.260 5.440 ;
        RECT  9.260 4.640 11.070 5.440 ;
        RECT  11.070 4.480 11.470 5.440 ;
        RECT  11.470 4.640 12.890 5.440 ;
        RECT  12.890 4.480 13.290 5.440 ;
        RECT  13.290 4.640 14.520 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.310 0.400 ;
        RECT  1.310 -0.400 1.710 0.560 ;
        RECT  1.710 -0.400 4.030 0.400 ;
        RECT  4.030 -0.400 4.040 1.020 ;
        RECT  4.040 -0.400 4.440 1.220 ;
        RECT  4.440 -0.400 4.450 1.020 ;
        RECT  4.450 -0.400 6.660 0.400 ;
        RECT  6.660 -0.400 7.060 1.410 ;
        RECT  7.060 -0.400 9.100 0.400 ;
        RECT  9.100 -0.400 9.500 1.390 ;
        RECT  9.500 -0.400 11.280 0.400 ;
        RECT  11.280 -0.400 11.290 0.790 ;
        RECT  11.290 -0.400 11.690 0.990 ;
        RECT  11.690 -0.400 11.700 0.790 ;
        RECT  11.700 -0.400 12.990 0.400 ;
        RECT  12.990 -0.400 13.390 0.560 ;
        RECT  13.390 -0.400 14.520 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  13.360 2.170 13.600 4.090 ;
        RECT  12.410 3.850 13.360 4.090 ;
        RECT  12.330 1.380 12.430 1.780 ;
        RECT  12.010 3.850 12.410 4.320 ;
        RECT  12.090 1.380 12.330 2.800 ;
        RECT  11.730 2.560 12.090 2.800 ;
        RECT  11.730 3.850 12.010 4.090 ;
        RECT  11.610 1.600 11.850 2.320 ;
        RECT  11.490 2.560 11.730 4.090 ;
        RECT  10.610 1.600 11.610 1.840 ;
        RECT  11.130 2.610 11.490 2.850 ;
        RECT  10.890 2.180 11.130 2.850 ;
        RECT  10.370 1.600 10.610 3.640 ;
        RECT  10.350 1.600 10.370 1.920 ;
        RECT  10.000 3.400 10.370 3.640 ;
        RECT  9.950 1.110 10.350 1.920 ;
        RECT  9.850 2.410 10.090 2.860 ;
        RECT  9.600 3.400 10.000 3.800 ;
        RECT  8.280 1.680 9.950 1.920 ;
        RECT  7.740 2.620 9.850 2.860 ;
        RECT  7.980 3.520 9.600 3.760 ;
        RECT  8.040 1.240 8.280 1.920 ;
        RECT  7.880 1.240 8.040 1.640 ;
        RECT  7.580 3.520 7.980 3.920 ;
        RECT  7.600 2.620 7.740 3.240 ;
        RECT  7.360 1.680 7.600 3.240 ;
        RECT  6.140 1.680 7.360 1.920 ;
        RECT  7.330 2.620 7.360 3.240 ;
        RECT  6.970 3.000 7.330 3.240 ;
        RECT  6.600 2.320 7.000 2.720 ;
        RECT  6.730 3.000 6.970 4.180 ;
        RECT  6.020 3.940 6.730 4.180 ;
        RECT  6.440 2.480 6.600 2.720 ;
        RECT  6.200 2.480 6.440 3.660 ;
        RECT  5.500 3.420 6.200 3.660 ;
        RECT  5.780 1.090 6.180 1.330 ;
        RECT  5.780 3.940 6.020 4.350 ;
        RECT  5.780 2.740 5.920 3.140 ;
        RECT  5.540 1.090 5.780 3.140 ;
        RECT  4.090 4.110 5.780 4.350 ;
        RECT  5.520 2.020 5.540 3.140 ;
        RECT  5.510 2.020 5.520 2.760 ;
        RECT  5.500 2.020 5.510 2.420 ;
        RECT  5.100 3.420 5.500 3.800 ;
        RECT  5.100 0.910 5.260 1.310 ;
        RECT  4.860 0.910 5.100 3.800 ;
        RECT  4.000 2.290 4.860 2.530 ;
        RECT  4.180 1.500 4.580 1.810 ;
        RECT  3.070 1.500 4.180 1.740 ;
        RECT  3.850 2.880 4.090 4.350 ;
        RECT  3.720 2.880 3.850 3.120 ;
        RECT  3.460 3.930 3.850 4.350 ;
        RECT  3.480 2.350 3.720 3.120 ;
        RECT  3.200 3.390 3.560 3.630 ;
        RECT  2.900 2.350 3.480 2.590 ;
        RECT  2.660 4.110 3.460 4.350 ;
        RECT  2.960 2.870 3.200 3.630 ;
        RECT  2.670 1.230 3.070 1.740 ;
        RECT  2.380 2.870 2.960 3.110 ;
        RECT  2.660 2.190 2.900 2.590 ;
        RECT  2.380 1.500 2.670 1.740 ;
        RECT  2.420 3.860 2.660 4.350 ;
        RECT  1.160 3.860 2.420 4.100 ;
        RECT  2.140 1.500 2.380 3.110 ;
        RECT  0.920 3.000 1.160 4.100 ;
        RECT  0.760 3.000 0.920 3.400 ;
        RECT  0.500 1.140 0.890 1.540 ;
        RECT  0.500 3.000 0.760 3.240 ;
        RECT  0.490 1.140 0.500 3.240 ;
        RECT  0.260 1.300 0.490 3.240 ;
    END
END DFFX2

MACRO DFFX1
    CLASS CORE ;
    FOREIGN DFFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ DFFXL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  11.180 3.570 11.380 3.810 ;
        RECT  11.380 1.540 11.390 3.810 ;
        RECT  11.390 1.160 11.670 3.810 ;
        RECT  11.670 2.390 11.680 2.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  9.620 3.050 10.010 3.450 ;
        RECT  10.010 3.050 10.100 3.740 ;
        RECT  9.870 0.690 10.270 1.100 ;
        RECT  10.100 3.050 10.360 3.770 ;
        RECT  10.360 3.050 10.450 3.740 ;
        RECT  10.450 3.050 10.820 3.290 ;
        RECT  10.270 0.860 10.820 1.100 ;
        RECT  10.820 0.860 11.060 3.290 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.270 1.780 1.930 ;
        RECT  1.780 1.280 1.830 1.930 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 1.030 2.650 ;
        RECT  1.030 2.380 1.430 2.780 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.510 5.440 ;
        RECT  1.510 4.480 1.910 5.440 ;
        RECT  1.910 4.640 6.490 5.440 ;
        RECT  6.490 4.480 6.890 5.440 ;
        RECT  6.890 4.640 8.800 5.440 ;
        RECT  8.800 4.480 9.200 5.440 ;
        RECT  9.200 4.640 10.420 5.440 ;
        RECT  10.420 4.480 10.820 5.440 ;
        RECT  10.820 4.640 11.880 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.360 0.400 ;
        RECT  1.360 -0.400 1.760 0.560 ;
        RECT  1.760 -0.400 4.030 0.400 ;
        RECT  4.030 -0.400 4.040 0.960 ;
        RECT  4.040 -0.400 4.440 1.160 ;
        RECT  4.440 -0.400 4.450 0.960 ;
        RECT  4.450 -0.400 6.660 0.400 ;
        RECT  6.660 -0.400 7.060 1.390 ;
        RECT  7.060 -0.400 9.100 0.400 ;
        RECT  9.100 -0.400 9.110 0.670 ;
        RECT  9.110 -0.400 9.510 0.870 ;
        RECT  9.510 -0.400 9.520 0.670 ;
        RECT  9.520 -0.400 10.700 0.400 ;
        RECT  10.700 -0.400 11.100 0.560 ;
        RECT  11.100 -0.400 11.880 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.300 1.430 10.540 2.770 ;
        RECT  9.930 1.430 10.300 1.670 ;
        RECT  9.060 2.530 10.300 2.770 ;
        RECT  9.740 4.050 10.020 4.290 ;
        RECT  9.610 2.000 9.780 2.240 ;
        RECT  9.500 3.940 9.740 4.290 ;
        RECT  9.370 1.600 9.610 2.240 ;
        RECT  9.050 3.940 9.500 4.180 ;
        RECT  8.280 1.600 9.370 1.840 ;
        RECT  9.050 2.130 9.060 2.770 ;
        RECT  8.810 2.130 9.050 4.180 ;
        RECT  8.660 2.130 8.810 2.530 ;
        RECT  7.600 0.760 8.610 1.000 ;
        RECT  8.270 1.290 8.280 1.840 ;
        RECT  8.030 1.290 8.270 4.370 ;
        RECT  7.880 1.290 8.030 1.690 ;
        RECT  7.770 3.970 8.030 4.370 ;
        RECT  7.600 2.310 7.640 2.710 ;
        RECT  7.440 0.760 7.600 2.710 ;
        RECT  7.360 0.760 7.440 4.180 ;
        RECT  6.140 1.680 7.360 1.920 ;
        RECT  7.200 2.390 7.360 4.180 ;
        RECT  6.210 3.940 7.200 4.180 ;
        RECT  6.680 2.320 6.920 3.660 ;
        RECT  5.690 3.420 6.680 3.660 ;
        RECT  5.970 3.940 6.210 4.370 ;
        RECT  5.780 0.850 6.180 1.250 ;
        RECT  4.120 4.130 5.970 4.370 ;
        RECT  5.760 2.740 5.920 3.140 ;
        RECT  5.760 1.010 5.780 1.250 ;
        RECT  5.520 1.010 5.760 3.140 ;
        RECT  5.450 3.420 5.690 3.850 ;
        RECT  5.500 1.490 5.520 1.890 ;
        RECT  4.860 3.610 5.450 3.850 ;
        RECT  5.220 0.760 5.240 1.160 ;
        RECT  5.000 0.760 5.220 2.390 ;
        RECT  4.980 0.840 5.000 2.390 ;
        RECT  4.860 2.150 4.980 2.390 ;
        RECT  4.600 2.150 4.860 3.850 ;
        RECT  4.240 2.150 4.600 2.560 ;
        RECT  4.180 1.430 4.580 1.830 ;
        RECT  3.920 2.150 4.240 2.550 ;
        RECT  3.100 1.590 4.180 1.830 ;
        RECT  3.880 2.890 4.120 4.370 ;
        RECT  2.880 2.890 3.880 3.130 ;
        RECT  3.480 3.940 3.880 4.370 ;
        RECT  2.360 3.420 3.560 3.660 ;
        RECT  1.080 3.940 3.480 4.180 ;
        RECT  2.940 0.910 3.100 1.830 ;
        RECT  2.700 0.910 2.940 2.050 ;
        RECT  2.640 2.330 2.880 3.130 ;
        RECT  2.360 1.810 2.700 2.050 ;
        RECT  2.120 1.810 2.360 3.660 ;
        RECT  0.840 3.450 1.080 4.180 ;
        RECT  0.530 0.860 0.880 1.260 ;
        RECT  0.680 3.450 0.840 3.850 ;
        RECT  0.530 3.450 0.680 3.690 ;
        RECT  0.480 0.860 0.530 3.690 ;
        RECT  0.290 0.980 0.480 3.690 ;
    END
END DFFX1

MACRO CLKINVXL
    CLASS CORE ;
    FOREIGN CLKINVXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 3.270 1.110 3.770 ;
        RECT  1.110 3.080 1.120 3.770 ;
        RECT  1.120 3.080 1.200 3.510 ;
        RECT  1.070 1.320 1.200 1.720 ;
        RECT  1.200 1.320 1.440 3.510 ;
        RECT  1.440 1.320 1.470 1.720 ;
        RECT  1.440 3.080 1.510 3.510 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.330 2.660 ;
        RECT  0.330 2.390 0.460 2.800 ;
        RECT  0.460 2.400 0.910 2.800 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.290 5.440 ;
        RECT  0.290 4.480 0.690 5.440 ;
        RECT  0.690 4.640 1.980 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.950 0.400 ;
        RECT  0.950 -0.400 1.350 0.560 ;
        RECT  1.350 -0.400 1.980 0.400 ;
        END
    END GND
END CLKINVXL

MACRO CLKINVX8
    CLASS CORE ;
    FOREIGN CLKINVX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKINVXL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.770 3.080 1.530 3.500 ;
        RECT  0.670 1.270 1.530 1.890 ;
        RECT  1.530 1.270 3.100 3.500 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.570 2.150 1.120 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.170 0.170 5.440 ;
        RECT  0.170 4.050 0.570 5.440 ;
        RECT  0.570 4.170 0.580 5.440 ;
        RECT  0.580 4.640 1.560 5.440 ;
        RECT  1.560 4.170 1.570 5.440 ;
        RECT  1.570 3.970 1.970 5.440 ;
        RECT  1.970 4.170 1.980 5.440 ;
        RECT  1.980 4.640 2.980 5.440 ;
        RECT  2.980 4.170 2.990 5.440 ;
        RECT  2.990 3.970 3.390 5.440 ;
        RECT  3.390 4.170 3.400 5.440 ;
        RECT  3.400 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.580 0.840 ;
        RECT  0.580 -0.400 1.510 0.400 ;
        RECT  1.510 -0.400 1.910 0.560 ;
        RECT  1.910 -0.400 4.620 0.400 ;
        END
    END GND
END CLKINVX8

MACRO CLKINVX4
    CLASS CORE ;
    FOREIGN CLKINVX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKINVXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.750 2.850 1.150 3.250 ;
        RECT  1.150 2.850 1.430 3.220 ;
        RECT  0.990 1.380 1.430 1.780 ;
        RECT  1.430 1.380 1.830 3.220 ;
        RECT  1.830 1.820 1.870 3.220 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.270 0.310 1.530 ;
        RECT  0.310 1.270 0.460 2.580 ;
        RECT  0.460 1.280 0.550 2.580 ;
        RECT  0.550 2.180 0.900 2.580 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.020 0.560 5.440 ;
        RECT  0.560 4.640 1.730 5.440 ;
        RECT  1.730 4.020 2.130 5.440 ;
        RECT  2.130 4.640 2.640 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.320 0.400 ;
        RECT  0.320 -0.400 0.720 0.560 ;
        RECT  0.720 -0.400 2.640 0.400 ;
        END
    END GND
END CLKINVX4

MACRO CLKINVX3
    CLASS CORE ;
    FOREIGN CLKINVX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKINVXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.770 2.930 0.910 3.780 ;
        RECT  0.910 2.930 1.310 3.910 ;
        RECT  1.310 2.930 1.370 3.170 ;
        RECT  1.290 0.900 1.370 1.800 ;
        RECT  1.370 0.900 1.610 3.170 ;
        RECT  1.610 0.900 1.690 1.960 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.210 2.650 ;
        RECT  0.210 1.840 0.450 2.650 ;
        RECT  0.450 2.040 0.460 2.650 ;
        RECT  0.460 2.040 1.070 2.440 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.250 5.440 ;
        RECT  0.250 2.950 0.490 5.440 ;
        RECT  0.490 4.640 1.730 5.440 ;
        RECT  1.730 4.480 2.130 5.440 ;
        RECT  2.130 4.640 2.640 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.460 0.400 ;
        RECT  0.460 -0.400 0.860 0.560 ;
        RECT  0.860 -0.400 2.640 0.400 ;
        END
    END GND
END CLKINVX3

MACRO CLKINVX2
    CLASS CORE ;
    FOREIGN CLKINVX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKINVXL ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.790 2.790 1.430 3.190 ;
        RECT  1.430 2.660 1.530 3.190 ;
        RECT  1.410 0.940 1.530 1.530 ;
        RECT  1.530 0.940 1.770 3.190 ;
        RECT  1.770 0.940 1.810 1.530 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.750 1.830 1.150 2.440 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.060 5.440 ;
        RECT  1.060 4.480 1.460 5.440 ;
        RECT  1.460 4.640 1.980 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.590 0.400 ;
        RECT  0.590 -0.400 0.990 1.540 ;
        RECT  0.990 -0.400 1.980 0.400 ;
        END
    END GND
END CLKINVX2

MACRO CLKINVX20
    CLASS CORE ;
    FOREIGN CLKINVX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKINVXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  7.030 2.800 11.130 3.820 ;
        RECT  11.130 2.500 11.430 3.820 ;
        RECT  6.370 1.230 11.430 1.870 ;
        RECT  11.430 1.200 12.990 3.840 ;
        RECT  12.990 1.200 13.090 3.820 ;
        RECT  13.090 1.260 13.250 3.820 ;
        RECT  13.250 1.260 13.530 2.790 ;
        RECT  13.530 1.390 14.180 2.790 ;
        RECT  14.180 1.680 14.330 2.790 ;
        RECT  14.330 1.680 14.730 3.720 ;
        RECT  14.730 1.680 14.840 2.790 ;
        RECT  14.840 1.690 15.490 2.790 ;
        RECT  15.490 1.680 15.850 2.790 ;
        RECT  15.850 1.680 16.250 3.720 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.010 2.020 1.520 2.420 ;
        RECT  1.520 1.830 1.780 2.420 ;
        RECT  1.780 2.020 1.910 2.420 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.250 5.440 ;
        RECT  0.250 2.740 0.650 5.440 ;
        RECT  0.650 4.640 1.980 5.440 ;
        RECT  1.980 4.190 1.990 5.440 ;
        RECT  1.990 3.990 2.390 5.440 ;
        RECT  2.390 4.190 2.400 5.440 ;
        RECT  2.400 4.640 3.470 5.440 ;
        RECT  3.470 4.210 3.480 5.440 ;
        RECT  3.480 4.010 3.880 5.440 ;
        RECT  3.880 4.210 3.890 5.440 ;
        RECT  3.890 4.640 5.000 5.440 ;
        RECT  5.000 4.350 5.010 5.440 ;
        RECT  5.010 4.150 5.410 5.440 ;
        RECT  5.410 4.350 5.420 5.440 ;
        RECT  5.420 4.640 6.310 5.440 ;
        RECT  6.310 3.580 6.710 5.440 ;
        RECT  6.710 4.640 7.750 5.440 ;
        RECT  7.750 4.130 8.150 5.440 ;
        RECT  8.150 4.640 9.190 5.440 ;
        RECT  9.190 4.130 9.590 5.440 ;
        RECT  9.590 4.640 10.630 5.440 ;
        RECT  10.630 4.130 11.030 5.440 ;
        RECT  11.030 4.640 12.070 5.440 ;
        RECT  12.070 4.130 12.470 5.440 ;
        RECT  12.470 4.640 13.610 5.440 ;
        RECT  13.610 3.080 14.010 5.440 ;
        RECT  14.010 4.640 15.130 5.440 ;
        RECT  15.130 3.080 15.530 5.440 ;
        RECT  15.530 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 2.050 0.400 ;
        RECT  2.050 -0.400 2.060 0.680 ;
        RECT  2.060 -0.400 2.460 0.880 ;
        RECT  2.460 -0.400 2.470 0.680 ;
        RECT  2.470 -0.400 3.720 0.400 ;
        RECT  3.720 -0.400 4.120 0.880 ;
        RECT  4.120 -0.400 5.470 0.400 ;
        RECT  5.470 -0.400 5.870 1.480 ;
        RECT  5.870 -0.400 7.200 0.400 ;
        RECT  7.200 -0.400 7.210 0.730 ;
        RECT  7.210 -0.400 7.610 0.930 ;
        RECT  7.610 -0.400 7.620 0.730 ;
        RECT  7.620 -0.400 8.530 0.400 ;
        RECT  8.530 -0.400 8.540 0.730 ;
        RECT  8.540 -0.400 8.940 0.930 ;
        RECT  8.940 -0.400 8.950 0.730 ;
        RECT  8.950 -0.400 9.880 0.400 ;
        RECT  9.880 -0.400 9.890 0.730 ;
        RECT  9.890 -0.400 10.290 0.930 ;
        RECT  10.290 -0.400 10.300 0.730 ;
        RECT  10.300 -0.400 11.160 0.400 ;
        RECT  11.160 -0.400 11.170 0.730 ;
        RECT  11.170 -0.400 11.570 0.930 ;
        RECT  11.570 -0.400 11.580 0.730 ;
        RECT  11.580 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.130 2.160 10.890 2.560 ;
        RECT  5.840 2.890 6.040 3.290 ;
        RECT  5.130 2.880 5.840 3.300 ;
        RECT  4.730 1.390 5.130 3.300 ;
        RECT  2.910 1.400 4.730 1.800 ;
        RECT  4.660 2.880 4.730 3.300 ;
        RECT  4.650 2.880 4.660 3.630 ;
        RECT  4.250 2.880 4.650 4.380 ;
        RECT  2.390 2.180 4.400 2.580 ;
        RECT  4.240 2.880 4.250 3.630 ;
        RECT  3.120 2.880 4.240 3.300 ;
        RECT  3.110 2.880 3.120 3.630 ;
        RECT  2.710 2.880 3.110 4.380 ;
        RECT  2.700 2.880 2.710 3.630 ;
        RECT  2.150 1.340 2.390 2.980 ;
        RECT  1.660 1.340 2.150 1.580 ;
        RECT  1.490 2.740 2.150 2.980 ;
        RECT  1.260 0.680 1.660 1.580 ;
        RECT  1.090 2.740 1.490 3.140 ;
    END
END CLKINVX20

MACRO CLKINVX1
    CLASS CORE ;
    FOREIGN CLKINVX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKINVXL ;
    SIZE 1.980 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.450 1.140 0.860 1.540 ;
        RECT  0.860 1.140 1.210 3.240 ;
        RECT  1.210 2.510 1.380 3.240 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.150 2.060 0.510 2.980 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.570 5.440 ;
        RECT  0.570 4.640 1.980 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.420 0.400 ;
        RECT  0.420 -0.400 0.820 0.560 ;
        RECT  0.820 -0.400 1.980 0.400 ;
        END
    END GND
END CLKINVX1

MACRO CLKINVX16
    CLASS CORE ;
    FOREIGN CLKINVX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKINVXL ;
    SIZE 14.520 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  5.600 2.840 10.510 3.840 ;
        RECT  10.510 2.510 10.770 3.840 ;
        RECT  5.860 1.200 10.770 1.880 ;
        RECT  10.770 1.200 12.330 3.840 ;
        RECT  12.330 2.500 13.700 3.840 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.690 2.180 0.770 2.580 ;
        RECT  0.770 2.180 0.860 2.640 ;
        RECT  0.860 2.180 1.090 2.650 ;
        RECT  1.090 2.390 1.120 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 3.350 0.180 5.440 ;
        RECT  0.180 3.150 0.580 5.440 ;
        RECT  0.580 3.350 0.590 5.440 ;
        RECT  0.590 4.640 1.760 5.440 ;
        RECT  1.760 4.080 1.770 5.440 ;
        RECT  1.770 3.600 2.170 5.440 ;
        RECT  2.170 4.080 2.180 5.440 ;
        RECT  2.180 4.640 3.300 5.440 ;
        RECT  3.300 4.080 3.310 5.440 ;
        RECT  3.310 3.600 3.710 5.440 ;
        RECT  3.710 4.080 3.720 5.440 ;
        RECT  3.720 4.640 4.850 5.440 ;
        RECT  4.850 4.370 4.860 5.440 ;
        RECT  4.860 4.170 5.260 5.440 ;
        RECT  5.260 4.370 5.270 5.440 ;
        RECT  5.270 4.640 6.320 5.440 ;
        RECT  6.320 4.360 6.330 5.440 ;
        RECT  6.330 4.160 6.730 5.440 ;
        RECT  6.730 4.360 6.740 5.440 ;
        RECT  6.740 4.640 7.930 5.440 ;
        RECT  7.930 4.360 7.940 5.440 ;
        RECT  7.940 4.160 8.340 5.440 ;
        RECT  8.340 4.360 8.350 5.440 ;
        RECT  8.350 4.640 9.430 5.440 ;
        RECT  9.430 4.360 9.440 5.440 ;
        RECT  9.440 4.160 9.840 5.440 ;
        RECT  9.840 4.360 9.850 5.440 ;
        RECT  9.850 4.640 10.950 5.440 ;
        RECT  10.950 4.360 10.960 5.440 ;
        RECT  10.960 4.160 11.360 5.440 ;
        RECT  11.360 4.360 11.370 5.440 ;
        RECT  11.370 4.640 12.520 5.440 ;
        RECT  12.520 4.360 12.530 5.440 ;
        RECT  12.530 4.160 12.930 5.440 ;
        RECT  12.930 4.360 12.940 5.440 ;
        RECT  12.940 4.640 13.930 5.440 ;
        RECT  13.930 4.360 13.940 5.440 ;
        RECT  13.940 4.160 14.340 5.440 ;
        RECT  14.340 4.360 14.350 5.440 ;
        RECT  14.350 4.640 14.520 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 2.120 0.400 ;
        RECT  2.120 -0.400 2.130 0.730 ;
        RECT  2.130 -0.400 2.530 0.930 ;
        RECT  2.530 -0.400 2.540 0.730 ;
        RECT  2.540 -0.400 3.380 0.400 ;
        RECT  3.380 -0.400 3.390 0.710 ;
        RECT  3.390 -0.400 3.790 0.910 ;
        RECT  3.790 -0.400 3.800 0.710 ;
        RECT  3.800 -0.400 5.250 0.400 ;
        RECT  5.250 -0.400 5.260 0.730 ;
        RECT  5.260 -0.400 5.660 0.850 ;
        RECT  5.660 -0.400 5.670 0.730 ;
        RECT  5.670 -0.400 6.640 0.400 ;
        RECT  6.640 -0.400 6.650 0.730 ;
        RECT  6.650 -0.400 7.050 0.930 ;
        RECT  7.050 -0.400 7.060 0.730 ;
        RECT  7.060 -0.400 8.000 0.400 ;
        RECT  8.000 -0.400 8.010 0.730 ;
        RECT  8.010 -0.400 8.410 0.930 ;
        RECT  8.410 -0.400 8.420 0.730 ;
        RECT  8.420 -0.400 9.340 0.400 ;
        RECT  9.340 -0.400 9.350 0.730 ;
        RECT  9.350 -0.400 9.750 0.930 ;
        RECT  9.750 -0.400 9.760 0.730 ;
        RECT  9.760 -0.400 14.520 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  7.710 2.160 10.080 2.560 ;
        RECT  5.070 2.150 7.710 2.570 ;
        RECT  4.650 1.380 5.070 3.230 ;
        RECT  2.980 1.380 4.650 1.800 ;
        RECT  4.490 2.810 4.650 3.230 ;
        RECT  4.480 2.810 4.490 3.320 ;
        RECT  4.080 2.810 4.480 3.800 ;
        RECT  1.730 2.070 4.300 2.470 ;
        RECT  4.070 2.810 4.080 3.320 ;
        RECT  2.940 2.810 4.070 3.230 ;
        RECT  2.780 1.390 2.980 1.790 ;
        RECT  2.930 2.810 2.940 3.320 ;
        RECT  2.530 2.810 2.930 3.800 ;
        RECT  2.520 2.810 2.530 3.320 ;
        RECT  1.490 1.370 1.730 3.190 ;
        RECT  1.330 1.370 1.490 1.770 ;
        RECT  1.340 2.950 1.490 3.190 ;
        RECT  0.940 2.950 1.340 3.350 ;
    END
END CLKINVX16

MACRO CLKINVX12
    CLASS CORE ;
    FOREIGN CLKINVX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKINVXL ;
    SIZE 12.540 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.730 2.880 9.450 3.840 ;
        RECT  4.640 1.200 9.450 1.880 ;
        RECT  9.450 1.200 11.010 3.840 ;
        RECT  11.010 1.200 11.020 1.860 ;
        RECT  11.010 2.520 11.310 3.840 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.770 1.280 0.860 2.480 ;
        RECT  0.860 1.270 1.010 2.480 ;
        RECT  1.010 1.270 1.120 1.530 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.940 5.440 ;
        RECT  0.940 4.340 0.950 5.440 ;
        RECT  0.950 4.140 1.350 5.440 ;
        RECT  1.350 4.340 1.360 5.440 ;
        RECT  1.360 4.640 2.480 5.440 ;
        RECT  2.480 4.480 2.880 5.440 ;
        RECT  2.880 4.640 4.050 5.440 ;
        RECT  4.050 4.480 4.450 5.440 ;
        RECT  4.450 4.640 5.480 5.440 ;
        RECT  5.480 4.320 5.490 5.440 ;
        RECT  5.490 4.120 5.890 5.440 ;
        RECT  5.890 4.320 5.900 5.440 ;
        RECT  5.900 4.640 7.050 5.440 ;
        RECT  7.050 4.360 7.060 5.440 ;
        RECT  7.060 4.160 7.460 5.440 ;
        RECT  7.460 4.360 7.470 5.440 ;
        RECT  7.470 4.640 8.510 5.440 ;
        RECT  8.510 4.360 8.520 5.440 ;
        RECT  8.520 4.160 8.920 5.440 ;
        RECT  8.920 4.360 8.930 5.440 ;
        RECT  8.930 4.640 10.170 5.440 ;
        RECT  10.170 4.360 10.180 5.440 ;
        RECT  10.180 4.160 10.580 5.440 ;
        RECT  10.580 4.360 10.590 5.440 ;
        RECT  10.590 4.640 11.530 5.440 ;
        RECT  11.530 4.360 11.540 5.440 ;
        RECT  11.540 4.160 11.940 5.440 ;
        RECT  11.940 4.360 11.950 5.440 ;
        RECT  11.950 4.640 12.540 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.240 0.400 ;
        RECT  1.240 -0.400 1.640 0.560 ;
        RECT  1.640 -0.400 3.390 0.400 ;
        RECT  3.390 -0.400 3.980 0.560 ;
        RECT  3.980 -0.400 4.220 1.800 ;
        RECT  4.220 -0.400 4.370 0.560 ;
        RECT  4.370 -0.400 5.280 0.400 ;
        RECT  5.280 -0.400 5.290 0.730 ;
        RECT  5.290 -0.400 5.690 0.930 ;
        RECT  5.690 -0.400 5.700 0.730 ;
        RECT  5.700 -0.400 6.640 0.400 ;
        RECT  6.640 -0.400 6.650 0.730 ;
        RECT  6.650 -0.400 7.050 0.930 ;
        RECT  7.050 -0.400 7.060 0.730 ;
        RECT  7.060 -0.400 12.540 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.390 2.160 9.130 2.560 ;
        RECT  3.670 2.210 4.390 2.510 ;
        RECT  3.590 2.210 3.670 3.800 ;
        RECT  3.350 1.550 3.590 3.800 ;
        RECT  2.450 1.550 3.350 1.790 ;
        RECT  3.270 2.840 3.350 3.800 ;
        RECT  2.180 3.330 3.270 3.630 ;
        RECT  1.640 2.070 2.900 2.470 ;
        RECT  2.050 0.840 2.450 1.800 ;
        RECT  1.780 3.280 2.180 3.680 ;
        RECT  1.400 2.070 1.640 3.030 ;
        RECT  0.560 2.790 1.400 3.030 ;
        RECT  0.490 2.790 0.560 3.190 ;
        RECT  0.250 1.390 0.490 3.190 ;
        RECT  0.160 2.790 0.250 3.190 ;
    END
END CLKINVX12

MACRO CLKBUFXL
    CLASS CORE ;
    FOREIGN CLKBUFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.950 1.530 3.210 ;
        RECT  1.530 2.930 2.170 3.330 ;
        RECT  2.070 1.400 2.170 1.800 ;
        RECT  2.170 1.400 2.410 3.330 ;
        RECT  2.410 1.400 2.470 1.960 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.740 2.150 0.820 2.550 ;
        RECT  0.820 2.150 0.860 2.640 ;
        RECT  0.860 2.150 1.120 2.650 ;
        RECT  1.120 2.150 1.140 2.550 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.150 5.440 ;
        RECT  1.150 4.480 1.550 5.440 ;
        RECT  1.550 4.640 2.640 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.060 0.400 ;
        RECT  1.060 -0.400 1.460 0.560 ;
        RECT  1.460 -0.400 2.640 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.720 2.070 1.880 2.470 ;
        RECT  1.480 1.550 1.720 2.470 ;
        RECT  0.570 1.550 1.480 1.790 ;
        RECT  0.460 2.930 0.630 3.330 ;
        RECT  0.460 1.390 0.570 1.790 ;
        RECT  0.230 1.390 0.460 3.330 ;
        RECT  0.220 1.390 0.230 3.250 ;
        RECT  0.170 1.390 0.220 1.790 ;
    END
END CLKBUFXL

MACRO CLKBUFX8
    CLASS CORE ;
    FOREIGN CLKBUFX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKBUFXL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.350 2.820 2.750 4.320 ;
        RECT  2.750 2.820 2.850 3.980 ;
        RECT  2.840 1.050 2.850 1.530 ;
        RECT  2.850 0.810 2.910 3.980 ;
        RECT  2.910 0.810 3.250 3.630 ;
        RECT  3.250 1.760 4.090 3.630 ;
        RECT  4.090 1.760 4.410 4.320 ;
        RECT  4.410 2.510 4.490 4.320 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.800 2.030 0.860 2.430 ;
        RECT  0.860 1.830 1.120 2.430 ;
        RECT  1.120 2.030 1.200 2.430 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.260 5.440 ;
        RECT  0.260 3.630 0.270 5.440 ;
        RECT  0.270 3.430 0.670 5.440 ;
        RECT  0.670 3.630 0.680 5.440 ;
        RECT  0.680 4.640 1.600 5.440 ;
        RECT  1.600 4.140 1.610 5.440 ;
        RECT  1.610 3.940 2.010 5.440 ;
        RECT  2.010 4.140 2.020 5.440 ;
        RECT  2.020 4.640 3.260 5.440 ;
        RECT  3.260 4.210 3.270 5.440 ;
        RECT  3.270 4.010 3.670 5.440 ;
        RECT  3.670 4.210 3.680 5.440 ;
        RECT  3.680 4.640 4.810 5.440 ;
        RECT  4.810 4.060 4.820 5.440 ;
        RECT  4.820 3.860 5.220 5.440 ;
        RECT  5.220 4.060 5.230 5.440 ;
        RECT  5.230 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 2.100 0.400 ;
        RECT  2.100 -0.400 2.110 0.670 ;
        RECT  2.110 -0.400 2.510 0.870 ;
        RECT  2.510 -0.400 2.520 0.670 ;
        RECT  2.520 -0.400 3.560 0.400 ;
        RECT  3.560 -0.400 3.570 0.670 ;
        RECT  3.570 -0.400 3.970 0.870 ;
        RECT  3.970 -0.400 3.980 0.670 ;
        RECT  3.980 -0.400 5.940 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.880 2.150 2.570 2.550 ;
        RECT  1.480 1.150 1.880 3.150 ;
        RECT  1.290 1.150 1.480 1.550 ;
        RECT  0.880 2.750 1.480 3.150 ;
    END
END CLKBUFX8

MACRO CLKBUFX4
    CLASS CORE ;
    FOREIGN CLKBUFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKBUFXL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.590 2.820 1.990 4.320 ;
        RECT  1.990 2.820 2.090 3.220 ;
        RECT  2.070 1.380 2.090 1.780 ;
        RECT  2.090 1.380 2.470 3.220 ;
        RECT  2.470 1.820 2.530 3.220 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 1.820 1.210 2.160 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.800 5.440 ;
        RECT  0.800 4.480 1.200 5.440 ;
        RECT  1.200 4.640 2.300 5.440 ;
        RECT  2.300 4.210 2.310 5.440 ;
        RECT  2.310 4.010 2.710 5.440 ;
        RECT  2.710 4.210 2.720 5.440 ;
        RECT  2.720 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.450 0.400 ;
        RECT  1.450 -0.400 1.460 0.740 ;
        RECT  1.460 -0.400 1.860 0.940 ;
        RECT  1.860 -0.400 1.870 0.740 ;
        RECT  1.870 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.690 2.150 1.850 2.550 ;
        RECT  1.450 1.310 1.690 2.550 ;
        RECT  0.570 1.310 1.450 1.550 ;
        RECT  0.410 1.260 0.570 1.550 ;
        RECT  0.410 2.750 0.570 3.150 ;
        RECT  0.170 1.260 0.410 3.150 ;
    END
END CLKBUFX4

MACRO CLKBUFX3
    CLASS CORE ;
    FOREIGN CLKBUFX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKBUFXL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 2.850 1.870 3.780 ;
        RECT  1.870 2.850 2.170 3.250 ;
        RECT  2.070 1.360 2.170 1.760 ;
        RECT  2.170 1.360 2.310 3.250 ;
        RECT  2.310 1.360 2.410 3.090 ;
        RECT  2.410 1.360 2.470 1.960 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 1.820 1.210 2.180 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.760 5.440 ;
        RECT  0.760 4.480 1.160 5.440 ;
        RECT  1.160 4.640 2.150 5.440 ;
        RECT  2.150 3.870 2.160 5.440 ;
        RECT  2.160 3.670 2.560 5.440 ;
        RECT  2.560 3.870 2.570 5.440 ;
        RECT  2.570 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.360 0.400 ;
        RECT  1.360 -0.400 1.370 0.830 ;
        RECT  1.370 -0.400 1.770 1.030 ;
        RECT  1.770 -0.400 1.780 0.830 ;
        RECT  1.780 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.720 2.150 1.880 2.550 ;
        RECT  1.480 1.310 1.720 2.550 ;
        RECT  0.570 1.310 1.480 1.550 ;
        RECT  0.410 1.260 0.570 1.550 ;
        RECT  0.410 2.750 0.570 3.150 ;
        RECT  0.170 1.260 0.410 3.150 ;
    END
END CLKBUFX3

MACRO CLKBUFX2
    CLASS CORE ;
    FOREIGN CLKBUFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKBUFXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.950 1.530 3.210 ;
        RECT  1.530 2.930 2.170 3.330 ;
        RECT  2.070 1.400 2.170 1.800 ;
        RECT  2.170 1.400 2.410 3.330 ;
        RECT  2.410 1.400 2.470 1.960 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.740 2.150 0.820 2.550 ;
        RECT  0.820 2.150 0.860 2.640 ;
        RECT  0.860 2.150 1.120 2.650 ;
        RECT  1.120 2.150 1.140 2.550 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.150 5.440 ;
        RECT  1.150 4.480 1.550 5.440 ;
        RECT  1.550 4.640 2.640 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.070 0.400 ;
        RECT  1.070 -0.400 1.470 0.560 ;
        RECT  1.470 -0.400 2.640 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.720 2.070 1.880 2.470 ;
        RECT  1.480 1.550 1.720 2.470 ;
        RECT  0.580 1.550 1.480 1.790 ;
        RECT  0.460 2.930 0.620 3.330 ;
        RECT  0.460 1.390 0.580 1.790 ;
        RECT  0.220 1.390 0.460 3.330 ;
        RECT  0.180 1.390 0.220 1.790 ;
    END
END CLKBUFX2

MACRO CLKBUFX20
    CLASS CORE ;
    FOREIGN CLKBUFX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKBUFXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  5.240 0.820 5.640 1.810 ;
        RECT  5.640 0.970 6.880 1.810 ;
        RECT  6.880 0.820 7.280 1.810 ;
        RECT  7.280 0.970 8.520 1.810 ;
        RECT  8.520 0.820 8.920 1.810 ;
        RECT  8.920 0.910 9.770 1.810 ;
        RECT  5.180 2.740 9.780 3.720 ;
        RECT  9.780 2.510 10.110 3.720 ;
        RECT  9.770 0.910 10.110 1.970 ;
        RECT  10.110 0.910 10.160 3.840 ;
        RECT  10.160 0.820 10.560 3.840 ;
        RECT  10.560 0.910 11.670 3.840 ;
        RECT  11.670 0.910 11.800 1.970 ;
        RECT  11.670 2.510 12.000 3.720 ;
        RECT  11.800 0.820 12.200 1.970 ;
        RECT  12.000 2.740 13.710 3.720 ;
        RECT  13.710 2.050 14.230 3.720 ;
        RECT  14.230 2.050 15.250 2.720 ;
        RECT  15.250 2.050 15.730 3.720 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.600 2.070 1.520 2.470 ;
        RECT  1.520 1.830 1.780 2.470 ;
        RECT  1.780 2.070 2.640 2.470 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 3.430 0.570 5.440 ;
        RECT  0.570 4.640 1.570 5.440 ;
        RECT  1.570 4.330 1.580 5.440 ;
        RECT  1.580 4.130 1.980 5.440 ;
        RECT  1.980 4.330 1.990 5.440 ;
        RECT  1.990 4.640 3.010 5.440 ;
        RECT  3.010 4.060 3.020 5.440 ;
        RECT  3.020 3.580 3.420 5.440 ;
        RECT  3.420 4.060 3.430 5.440 ;
        RECT  3.430 4.640 4.450 5.440 ;
        RECT  4.450 3.790 4.460 5.440 ;
        RECT  4.460 3.040 4.860 5.440 ;
        RECT  4.860 3.790 4.870 5.440 ;
        RECT  4.870 4.640 5.890 5.440 ;
        RECT  5.890 4.230 5.900 5.440 ;
        RECT  5.900 4.030 6.300 5.440 ;
        RECT  6.300 4.230 6.310 5.440 ;
        RECT  6.310 4.640 7.330 5.440 ;
        RECT  7.330 4.230 7.340 5.440 ;
        RECT  7.340 4.030 7.740 5.440 ;
        RECT  7.740 4.230 7.750 5.440 ;
        RECT  7.750 4.640 8.770 5.440 ;
        RECT  8.770 4.310 8.780 5.440 ;
        RECT  8.780 4.110 9.180 5.440 ;
        RECT  9.180 4.310 9.190 5.440 ;
        RECT  9.190 4.640 10.210 5.440 ;
        RECT  10.210 4.320 10.220 5.440 ;
        RECT  10.220 4.120 10.620 5.440 ;
        RECT  10.620 4.320 10.630 5.440 ;
        RECT  10.630 4.640 11.650 5.440 ;
        RECT  11.650 4.330 11.660 5.440 ;
        RECT  11.660 4.130 12.060 5.440 ;
        RECT  12.060 4.330 12.070 5.440 ;
        RECT  12.070 4.640 13.090 5.440 ;
        RECT  13.090 4.230 13.100 5.440 ;
        RECT  13.100 4.030 13.500 5.440 ;
        RECT  13.500 4.230 13.510 5.440 ;
        RECT  13.510 4.640 14.530 5.440 ;
        RECT  14.530 3.790 14.540 5.440 ;
        RECT  14.540 3.040 14.940 5.440 ;
        RECT  14.940 3.790 14.950 5.440 ;
        RECT  14.950 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 2.900 0.400 ;
        RECT  2.900 -0.400 3.300 0.560 ;
        RECT  3.300 -0.400 4.470 0.400 ;
        RECT  4.470 -0.400 4.480 1.270 ;
        RECT  4.480 -0.400 4.880 1.760 ;
        RECT  4.880 -0.400 4.890 1.270 ;
        RECT  4.890 -0.400 6.060 0.400 ;
        RECT  6.060 -0.400 6.460 0.560 ;
        RECT  6.460 -0.400 7.700 0.400 ;
        RECT  7.700 -0.400 8.100 0.560 ;
        RECT  8.100 -0.400 9.340 0.400 ;
        RECT  9.340 -0.400 9.740 0.560 ;
        RECT  9.740 -0.400 10.980 0.400 ;
        RECT  10.980 -0.400 11.380 0.560 ;
        RECT  11.380 -0.400 12.550 0.400 ;
        RECT  12.550 -0.400 12.560 1.220 ;
        RECT  12.560 -0.400 12.960 1.710 ;
        RECT  12.960 -0.400 12.970 1.220 ;
        RECT  12.970 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.120 2.070 9.190 2.470 ;
        RECT  4.120 2.750 4.140 4.250 ;
        RECT  3.740 0.800 4.120 4.250 ;
        RECT  3.720 0.800 3.740 3.150 ;
        RECT  2.280 1.080 3.720 1.500 ;
        RECT  2.710 2.750 3.720 3.150 ;
        RECT  2.700 2.740 2.710 3.240 ;
        RECT  2.300 2.740 2.700 3.720 ;
        RECT  2.290 2.740 2.300 3.240 ;
        RECT  1.080 2.740 2.290 3.160 ;
        RECT  2.080 1.090 2.280 1.490 ;
        RECT  0.880 2.750 1.080 3.150 ;
    END
END CLKBUFX20

MACRO CLKBUFX1
    CLASS CORE ;
    FOREIGN CLKBUFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKBUFXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.950 1.530 3.210 ;
        RECT  1.530 2.930 2.170 3.330 ;
        RECT  2.070 1.400 2.170 1.830 ;
        RECT  2.170 1.400 2.410 3.330 ;
        RECT  2.410 1.400 2.470 1.960 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.740 2.150 0.820 2.550 ;
        RECT  0.820 2.150 0.860 2.640 ;
        RECT  0.860 2.150 1.120 2.650 ;
        RECT  1.120 2.150 1.140 2.550 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.150 5.440 ;
        RECT  1.150 4.480 1.550 5.440 ;
        RECT  1.550 4.640 2.640 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.060 0.400 ;
        RECT  1.060 -0.400 1.460 0.560 ;
        RECT  1.460 -0.400 2.640 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.720 2.070 1.880 2.470 ;
        RECT  1.480 1.470 1.720 2.470 ;
        RECT  0.570 1.470 1.480 1.710 ;
        RECT  0.460 2.930 0.620 3.330 ;
        RECT  0.460 1.390 0.570 1.790 ;
        RECT  0.220 1.390 0.460 3.330 ;
        RECT  0.170 1.390 0.220 1.790 ;
    END
END CLKBUFX1

MACRO CLKBUFX16
    CLASS CORE ;
    FOREIGN CLKBUFX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKBUFXL ;
    SIZE 13.860 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.520 0.820 4.920 1.800 ;
        RECT  4.920 0.970 5.910 1.800 ;
        RECT  5.910 0.820 6.560 1.800 ;
        RECT  6.560 0.970 7.790 1.800 ;
        RECT  4.480 2.740 7.800 3.740 ;
        RECT  7.790 0.970 7.800 1.960 ;
        RECT  7.800 2.520 8.130 3.740 ;
        RECT  7.800 0.820 8.130 1.960 ;
        RECT  8.130 0.820 8.200 3.840 ;
        RECT  8.200 0.910 9.440 3.840 ;
        RECT  9.440 0.820 9.690 3.840 ;
        RECT  9.690 0.820 9.840 1.950 ;
        RECT  9.840 1.170 9.850 1.950 ;
        RECT  9.690 2.530 10.020 3.740 ;
        RECT  10.020 2.740 13.540 3.740 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.680 2.030 1.520 2.430 ;
        RECT  1.520 1.830 1.780 2.430 ;
        RECT  1.780 2.030 2.720 2.430 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.880 5.440 ;
        RECT  0.880 3.870 0.890 5.440 ;
        RECT  0.890 3.670 1.290 5.440 ;
        RECT  1.290 3.870 1.300 5.440 ;
        RECT  1.300 4.640 2.320 5.440 ;
        RECT  2.320 3.900 2.330 5.440 ;
        RECT  2.330 3.700 2.730 5.440 ;
        RECT  2.730 3.900 2.740 5.440 ;
        RECT  2.740 4.640 3.760 5.440 ;
        RECT  3.760 3.640 3.770 5.440 ;
        RECT  3.770 2.890 4.170 5.440 ;
        RECT  4.170 3.640 4.180 5.440 ;
        RECT  4.180 4.640 5.200 5.440 ;
        RECT  5.200 4.330 5.210 5.440 ;
        RECT  5.210 4.130 5.610 5.440 ;
        RECT  5.610 4.330 5.620 5.440 ;
        RECT  5.620 4.640 6.640 5.440 ;
        RECT  6.640 4.330 6.650 5.440 ;
        RECT  6.650 4.130 7.050 5.440 ;
        RECT  7.050 4.330 7.060 5.440 ;
        RECT  7.060 4.640 8.080 5.440 ;
        RECT  8.080 4.270 8.090 5.440 ;
        RECT  8.090 4.150 8.490 5.440 ;
        RECT  8.490 4.270 8.500 5.440 ;
        RECT  8.500 4.640 9.520 5.440 ;
        RECT  9.520 4.330 9.530 5.440 ;
        RECT  9.530 4.210 9.930 5.440 ;
        RECT  9.930 4.330 9.940 5.440 ;
        RECT  9.940 4.640 10.960 5.440 ;
        RECT  10.960 4.230 10.970 5.440 ;
        RECT  10.970 4.030 11.370 5.440 ;
        RECT  11.370 4.230 11.380 5.440 ;
        RECT  11.380 4.640 12.400 5.440 ;
        RECT  12.400 4.230 12.410 5.440 ;
        RECT  12.410 4.030 12.810 5.440 ;
        RECT  12.810 4.230 12.820 5.440 ;
        RECT  12.820 4.640 13.860 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 2.180 0.400 ;
        RECT  2.180 -0.400 2.580 0.560 ;
        RECT  2.580 -0.400 3.750 0.400 ;
        RECT  3.750 -0.400 3.760 1.270 ;
        RECT  3.760 -0.400 4.160 1.760 ;
        RECT  4.160 -0.400 4.170 1.270 ;
        RECT  4.170 -0.400 5.340 0.400 ;
        RECT  5.340 -0.400 5.740 0.560 ;
        RECT  5.740 -0.400 6.980 0.400 ;
        RECT  6.980 -0.400 7.380 0.560 ;
        RECT  7.380 -0.400 8.620 0.400 ;
        RECT  8.620 -0.400 9.020 0.560 ;
        RECT  9.020 -0.400 10.190 0.400 ;
        RECT  10.190 -0.400 10.200 1.220 ;
        RECT  10.200 -0.400 10.600 1.710 ;
        RECT  10.600 -0.400 10.610 1.220 ;
        RECT  10.610 -0.400 13.860 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.820 2.070 7.380 2.470 ;
        RECT  3.460 2.060 5.820 2.480 ;
        RECT  3.450 2.060 3.460 3.520 ;
        RECT  3.410 2.060 3.450 4.270 ;
        RECT  3.400 1.290 3.410 4.270 ;
        RECT  3.050 0.800 3.400 4.270 ;
        RECT  3.040 0.800 3.050 3.520 ;
        RECT  3.000 0.800 3.040 2.480 ;
        RECT  2.020 2.750 3.040 3.170 ;
        RECT  2.990 1.080 3.000 2.480 ;
        RECT  1.560 1.080 2.990 1.500 ;
        RECT  2.010 2.750 2.020 3.230 ;
        RECT  1.610 2.750 2.010 3.710 ;
        RECT  1.600 2.750 1.610 3.230 ;
        RECT  0.580 2.750 1.600 3.170 ;
        RECT  1.360 1.090 1.560 1.490 ;
        RECT  0.570 2.750 0.580 3.230 ;
        RECT  0.170 2.750 0.570 3.710 ;
        RECT  0.160 2.750 0.170 3.230 ;
    END
END CLKBUFX16

MACRO CLKBUFX12
    CLASS CORE ;
    FOREIGN CLKBUFX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ CLKBUFXL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.250 0.820 4.650 1.800 ;
        RECT  4.650 0.970 5.890 1.800 ;
        RECT  5.890 0.820 6.290 1.800 ;
        RECT  6.290 0.970 7.530 1.800 ;
        RECT  7.530 0.820 7.790 1.800 ;
        RECT  3.830 2.740 7.800 3.740 ;
        RECT  7.790 0.820 7.930 1.950 ;
        RECT  7.800 2.520 8.130 3.740 ;
        RECT  7.930 0.970 8.130 1.950 ;
        RECT  8.130 0.970 9.690 3.740 ;
        RECT  9.690 0.970 9.700 1.950 ;
        RECT  9.690 2.650 10.450 3.740 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.710 2.030 0.860 2.430 ;
        RECT  0.860 1.830 1.120 2.430 ;
        RECT  1.120 2.030 2.250 2.430 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.360 5.440 ;
        RECT  0.360 3.920 0.370 5.440 ;
        RECT  0.370 3.720 0.770 5.440 ;
        RECT  0.770 3.920 0.780 5.440 ;
        RECT  0.780 4.640 1.630 5.440 ;
        RECT  1.630 3.920 1.640 5.440 ;
        RECT  1.640 3.720 2.040 5.440 ;
        RECT  2.040 3.920 2.050 5.440 ;
        RECT  2.050 4.640 3.020 5.440 ;
        RECT  3.020 3.960 3.030 5.440 ;
        RECT  3.030 3.480 3.430 5.440 ;
        RECT  3.430 3.960 3.440 5.440 ;
        RECT  3.440 4.640 4.550 5.440 ;
        RECT  4.550 4.230 4.560 5.440 ;
        RECT  4.560 4.030 4.960 5.440 ;
        RECT  4.960 4.230 4.970 5.440 ;
        RECT  4.970 4.640 6.140 5.440 ;
        RECT  6.140 4.230 6.150 5.440 ;
        RECT  6.150 4.030 6.550 5.440 ;
        RECT  6.550 4.230 6.560 5.440 ;
        RECT  6.560 4.640 7.690 5.440 ;
        RECT  7.690 4.230 7.700 5.440 ;
        RECT  7.700 4.030 8.100 5.440 ;
        RECT  8.100 4.230 8.110 5.440 ;
        RECT  8.110 4.640 9.210 5.440 ;
        RECT  9.210 4.230 9.220 5.440 ;
        RECT  9.220 4.030 9.620 5.440 ;
        RECT  9.620 4.230 9.630 5.440 ;
        RECT  9.630 4.640 10.640 5.440 ;
        RECT  10.640 4.230 10.650 5.440 ;
        RECT  10.650 4.030 11.050 5.440 ;
        RECT  11.050 4.230 11.060 5.440 ;
        RECT  11.060 4.640 11.220 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.960 0.400 ;
        RECT  1.960 -0.400 1.970 1.220 ;
        RECT  1.970 -0.400 2.370 1.710 ;
        RECT  2.370 -0.400 2.380 1.220 ;
        RECT  2.380 -0.400 3.480 0.400 ;
        RECT  3.480 -0.400 3.490 1.130 ;
        RECT  3.490 -0.400 3.890 1.620 ;
        RECT  3.890 -0.400 3.900 1.130 ;
        RECT  3.900 -0.400 5.070 0.400 ;
        RECT  5.070 -0.400 5.470 0.560 ;
        RECT  5.470 -0.400 6.710 0.400 ;
        RECT  6.710 -0.400 7.110 0.560 ;
        RECT  7.110 -0.400 8.350 0.400 ;
        RECT  8.350 -0.400 8.750 0.560 ;
        RECT  8.750 -0.400 11.220 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.510 2.070 7.340 2.470 ;
        RECT  3.140 2.060 5.510 2.480 ;
        RECT  3.130 1.220 3.140 3.160 ;
        RECT  2.730 0.730 3.130 3.160 ;
        RECT  2.720 1.220 2.730 3.160 ;
        RECT  1.190 2.740 2.720 3.160 ;
        RECT  0.990 2.750 1.190 3.150 ;
    END
END CLKBUFX12

MACRO BUFXL
    CLASS CORE ;
    FOREIGN BUFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.270 1.630 1.530 ;
        RECT  1.630 1.260 2.050 1.540 ;
        RECT  2.030 2.840 2.190 3.240 ;
        RECT  2.190 2.640 2.210 3.240 ;
        RECT  2.050 1.150 2.210 1.550 ;
        RECT  2.210 1.150 2.450 3.240 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.770 1.790 1.210 2.360 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.150 5.440 ;
        RECT  1.150 4.480 1.550 5.440 ;
        RECT  1.550 4.640 2.640 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.130 0.400 ;
        RECT  1.130 -0.400 1.530 0.560 ;
        RECT  1.530 -0.400 2.640 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.730 1.830 1.910 2.230 ;
        RECT  1.490 1.830 1.730 3.010 ;
        RECT  0.610 2.770 1.490 3.010 ;
        RECT  0.450 1.150 0.610 1.550 ;
        RECT  0.450 2.770 0.610 3.170 ;
        RECT  0.210 1.150 0.450 3.170 ;
    END
END BUFXL

MACRO BUFX8
    CLASS CORE ;
    FOREIGN BUFX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BUFXL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.320 2.840 2.850 3.240 ;
        RECT  2.250 1.390 2.850 1.790 ;
        RECT  2.850 1.390 3.990 3.280 ;
        RECT  3.990 1.760 4.410 3.280 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.560 2.180 0.860 2.580 ;
        RECT  0.860 2.180 0.960 2.650 ;
        RECT  0.960 2.260 1.110 2.650 ;
        RECT  1.110 2.390 1.120 2.650 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.740 0.560 5.440 ;
        RECT  0.560 4.640 1.610 5.440 ;
        RECT  1.610 4.100 2.010 5.440 ;
        RECT  2.010 4.640 3.080 5.440 ;
        RECT  3.080 4.300 3.090 5.440 ;
        RECT  3.090 4.100 3.490 5.440 ;
        RECT  3.490 4.300 3.500 5.440 ;
        RECT  3.500 4.640 4.470 5.440 ;
        RECT  4.470 4.300 4.480 5.440 ;
        RECT  4.480 4.100 4.880 5.440 ;
        RECT  4.880 4.300 4.890 5.440 ;
        RECT  4.890 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.560 0.560 ;
        RECT  0.560 -0.400 1.600 0.400 ;
        RECT  1.600 -0.400 1.610 0.910 ;
        RECT  1.610 -0.400 2.010 1.110 ;
        RECT  2.010 -0.400 2.020 0.910 ;
        RECT  2.020 -0.400 2.910 0.400 ;
        RECT  2.910 -0.400 2.920 0.910 ;
        RECT  2.920 -0.400 3.320 1.110 ;
        RECT  3.320 -0.400 3.330 0.910 ;
        RECT  3.330 -0.400 4.200 0.400 ;
        RECT  4.200 -0.400 4.210 0.910 ;
        RECT  4.210 -0.400 4.610 1.110 ;
        RECT  4.610 -0.400 4.620 0.910 ;
        RECT  4.620 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.370 2.130 2.570 2.530 ;
        RECT  1.910 2.120 2.370 2.540 ;
        RECT  1.900 1.380 1.910 2.540 ;
        RECT  1.500 1.380 1.900 3.330 ;
        RECT  1.490 1.380 1.500 2.540 ;
        RECT  0.780 2.930 1.500 3.330 ;
        RECT  0.910 1.380 1.490 1.800 ;
        RECT  0.710 1.390 0.910 1.790 ;
    END
END BUFX8

MACRO BUFX4
    CLASS CORE ;
    FOREIGN BUFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BUFXL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.760 3.210 2.090 4.190 ;
        RECT  1.700 0.820 2.090 1.800 ;
        RECT  2.090 0.820 2.100 4.190 ;
        RECT  2.100 1.170 2.110 4.190 ;
        RECT  2.110 1.520 2.370 4.190 ;
        RECT  2.370 2.380 2.530 4.190 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.690 1.990 0.700 2.270 ;
        RECT  0.700 1.990 0.860 2.420 ;
        RECT  0.860 1.830 1.100 2.420 ;
        RECT  1.100 1.830 1.120 2.270 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 3.700 1.000 5.440 ;
        RECT  1.000 3.210 1.400 5.440 ;
        RECT  1.400 3.700 1.410 5.440 ;
        RECT  1.410 4.640 2.730 5.440 ;
        RECT  2.730 4.480 3.130 5.440 ;
        RECT  3.130 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.930 0.400 ;
        RECT  0.930 -0.400 0.940 1.220 ;
        RECT  0.940 -0.400 1.340 1.420 ;
        RECT  1.340 -0.400 1.350 1.220 ;
        RECT  1.350 -0.400 2.450 0.400 ;
        RECT  2.450 -0.400 2.460 1.040 ;
        RECT  2.460 -0.400 2.860 1.240 ;
        RECT  2.860 -0.400 2.870 1.040 ;
        RECT  2.870 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.610 2.070 1.850 2.940 ;
        RECT  0.580 2.700 1.610 2.940 ;
        RECT  0.420 1.080 0.580 1.480 ;
        RECT  0.420 2.700 0.580 3.820 ;
        RECT  0.180 1.080 0.420 3.820 ;
    END
END BUFX4

MACRO BUFX3
    CLASS CORE ;
    FOREIGN BUFX3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BUFXL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.700 1.060 1.830 1.460 ;
        RECT  1.760 3.080 2.090 4.100 ;
        RECT  1.830 1.060 2.090 1.800 ;
        RECT  2.090 1.060 2.100 4.100 ;
        RECT  2.100 1.120 2.110 4.100 ;
        RECT  2.110 1.520 2.370 4.100 ;
        RECT  2.370 2.940 2.530 4.100 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.690 1.820 0.700 2.100 ;
        RECT  0.700 1.820 1.110 2.250 ;
        RECT  1.110 1.820 1.120 2.100 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 3.610 1.000 5.440 ;
        RECT  1.000 3.120 1.400 5.440 ;
        RECT  1.400 3.610 1.410 5.440 ;
        RECT  1.410 4.640 2.730 5.440 ;
        RECT  2.730 4.480 3.130 5.440 ;
        RECT  3.130 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.930 0.400 ;
        RECT  0.930 -0.400 0.940 1.220 ;
        RECT  0.940 -0.400 1.340 1.420 ;
        RECT  1.340 -0.400 1.350 1.220 ;
        RECT  1.350 -0.400 2.450 0.400 ;
        RECT  2.450 -0.400 2.460 1.040 ;
        RECT  2.460 -0.400 2.860 1.240 ;
        RECT  2.860 -0.400 2.870 1.040 ;
        RECT  2.870 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.610 2.070 1.850 2.800 ;
        RECT  0.580 2.560 1.610 2.800 ;
        RECT  0.420 1.080 0.580 1.480 ;
        RECT  0.420 2.560 0.580 3.820 ;
        RECT  0.180 1.080 0.420 3.820 ;
    END
END BUFX3

MACRO BUFX2
    CLASS CORE ;
    FOREIGN BUFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BUFXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.270 1.630 1.530 ;
        RECT  1.630 1.260 2.070 1.540 ;
        RECT  2.070 2.800 2.190 3.200 ;
        RECT  2.190 2.640 2.230 3.200 ;
        RECT  2.070 0.930 2.230 1.540 ;
        RECT  2.230 0.930 2.470 3.200 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.770 1.820 1.210 2.240 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.160 5.440 ;
        RECT  1.160 4.480 1.560 5.440 ;
        RECT  1.560 4.640 2.640 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.170 0.400 ;
        RECT  1.170 -0.400 1.570 0.560 ;
        RECT  1.570 -0.400 2.640 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.790 2.010 1.920 2.410 ;
        RECT  1.550 2.010 1.790 3.000 ;
        RECT  1.520 2.010 1.550 2.410 ;
        RECT  0.660 2.760 1.550 3.000 ;
        RECT  0.500 1.150 0.660 1.550 ;
        RECT  0.500 2.760 0.660 3.180 ;
        RECT  0.260 1.150 0.500 3.180 ;
    END
END BUFX2

MACRO BUFX20
    CLASS CORE ;
    FOREIGN BUFX20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BUFXL ;
    SIZE 11.880 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.330 2.840 4.730 3.820 ;
        RECT  4.730 2.940 4.950 3.820 ;
        RECT  4.950 2.940 5.600 3.620 ;
        RECT  5.600 2.940 5.880 3.820 ;
        RECT  5.880 2.840 6.280 3.820 ;
        RECT  6.280 2.940 7.280 3.620 ;
        RECT  7.280 2.520 7.420 3.620 ;
        RECT  7.420 2.520 7.470 3.820 ;
        RECT  4.330 1.200 7.470 1.880 ;
        RECT  7.470 1.200 9.030 3.840 ;
        RECT  9.030 2.510 9.350 3.820 ;
        RECT  9.350 2.940 9.570 3.820 ;
        RECT  9.570 2.940 10.230 3.620 ;
        RECT  9.030 1.200 10.320 1.880 ;
        RECT  10.230 2.940 10.470 3.820 ;
        RECT  10.470 2.840 10.870 3.820 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.070 2.180 2.470 ;
        RECT  2.180 2.070 2.440 2.650 ;
        RECT  2.440 2.070 3.020 2.470 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.420 5.440 ;
        RECT  0.420 4.010 0.820 5.440 ;
        RECT  0.820 4.640 1.840 5.440 ;
        RECT  1.840 4.210 1.850 5.440 ;
        RECT  1.850 4.010 2.250 5.440 ;
        RECT  2.250 4.210 2.260 5.440 ;
        RECT  2.260 4.640 3.680 5.440 ;
        RECT  3.680 4.330 3.690 5.440 ;
        RECT  3.690 4.130 4.090 5.440 ;
        RECT  4.090 4.330 4.100 5.440 ;
        RECT  4.100 4.640 5.100 5.440 ;
        RECT  5.100 4.480 5.500 5.440 ;
        RECT  5.500 4.640 6.640 5.440 ;
        RECT  6.640 4.330 6.650 5.440 ;
        RECT  6.650 4.130 7.050 5.440 ;
        RECT  7.050 4.330 7.060 5.440 ;
        RECT  7.060 4.640 8.180 5.440 ;
        RECT  8.180 4.480 8.580 5.440 ;
        RECT  8.580 4.640 9.720 5.440 ;
        RECT  9.720 4.330 9.730 5.440 ;
        RECT  9.730 4.130 10.130 5.440 ;
        RECT  10.130 4.330 10.140 5.440 ;
        RECT  10.140 4.640 11.260 5.440 ;
        RECT  11.260 3.170 11.270 5.440 ;
        RECT  11.270 2.970 11.670 5.440 ;
        RECT  11.670 3.170 11.680 5.440 ;
        RECT  11.680 4.640 11.880 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.020 0.400 ;
        RECT  1.020 -0.400 1.030 0.910 ;
        RECT  1.030 -0.400 1.430 1.110 ;
        RECT  1.430 -0.400 1.440 0.910 ;
        RECT  1.440 -0.400 2.310 0.400 ;
        RECT  2.310 -0.400 2.320 0.910 ;
        RECT  2.320 -0.400 2.720 1.110 ;
        RECT  2.720 -0.400 2.730 0.910 ;
        RECT  2.730 -0.400 3.690 0.400 ;
        RECT  3.690 -0.400 4.090 0.920 ;
        RECT  4.090 -0.400 5.000 0.400 ;
        RECT  5.000 -0.400 5.010 0.730 ;
        RECT  5.010 -0.400 5.410 0.930 ;
        RECT  5.410 -0.400 5.420 0.730 ;
        RECT  5.420 -0.400 6.340 0.400 ;
        RECT  6.340 -0.400 6.350 0.730 ;
        RECT  6.350 -0.400 6.750 0.930 ;
        RECT  6.750 -0.400 6.760 0.730 ;
        RECT  6.760 -0.400 7.680 0.400 ;
        RECT  7.680 -0.400 7.690 0.730 ;
        RECT  7.690 -0.400 8.090 0.930 ;
        RECT  8.090 -0.400 8.100 0.730 ;
        RECT  8.100 -0.400 8.970 0.400 ;
        RECT  8.970 -0.400 8.980 0.730 ;
        RECT  8.980 -0.400 9.380 0.930 ;
        RECT  9.380 -0.400 9.390 0.730 ;
        RECT  9.390 -0.400 11.880 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.660 2.160 6.990 2.560 ;
        RECT  3.700 2.150 5.660 2.570 ;
        RECT  3.280 1.380 3.700 3.340 ;
        RECT  1.850 1.380 3.280 1.800 ;
        RECT  1.250 2.920 3.280 3.340 ;
        RECT  1.650 1.390 1.850 1.790 ;
        RECT  1.050 2.930 1.250 3.330 ;
    END
END BUFX20

MACRO BUFX1
    CLASS CORE ;
    FOREIGN BUFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BUFXL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.040 2.790 2.090 3.190 ;
        RECT  2.000 1.010 2.180 1.410 ;
        RECT  2.090 2.660 2.190 3.190 ;
        RECT  2.190 2.640 2.200 3.190 ;
        RECT  2.180 1.010 2.200 1.530 ;
        RECT  2.200 1.010 2.430 3.190 ;
        RECT  2.430 1.270 2.440 3.190 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.500 1.760 0.900 2.160 ;
        RECT  0.900 1.830 1.120 2.090 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.120 5.440 ;
        RECT  1.120 4.480 1.520 5.440 ;
        RECT  1.520 4.640 2.640 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.120 0.400 ;
        RECT  1.120 -0.400 1.520 0.560 ;
        RECT  1.520 -0.400 2.640 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.720 1.760 1.810 2.160 ;
        RECT  1.480 1.160 1.720 3.070 ;
        RECT  0.610 1.160 1.480 1.400 ;
        RECT  0.590 2.830 1.480 3.070 ;
        RECT  0.210 1.080 0.610 1.480 ;
        RECT  0.190 2.750 0.590 3.150 ;
    END
END BUFX1

MACRO BUFX16
    CLASS CORE ;
    FOREIGN BUFX16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BUFXL ;
    SIZE 9.240 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.190 2.840 3.200 3.520 ;
        RECT  3.200 2.840 3.600 3.820 ;
        RECT  3.600 2.840 4.740 3.520 ;
        RECT  4.740 2.840 5.140 3.820 ;
        RECT  5.140 2.840 6.280 3.520 ;
        RECT  6.280 2.840 6.710 3.840 ;
        RECT  6.710 2.500 6.810 3.840 ;
        RECT  3.330 1.200 6.810 1.880 ;
        RECT  6.810 1.200 8.370 3.840 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.750 2.070 1.520 2.470 ;
        RECT  1.520 2.070 1.780 2.650 ;
        RECT  1.780 2.070 2.250 2.470 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.880 5.440 ;
        RECT  0.880 4.080 0.890 5.440 ;
        RECT  0.890 3.600 1.290 5.440 ;
        RECT  1.290 4.080 1.300 5.440 ;
        RECT  1.300 4.640 2.420 5.440 ;
        RECT  2.420 3.990 2.430 5.440 ;
        RECT  2.430 3.790 2.830 5.440 ;
        RECT  2.830 3.990 2.840 5.440 ;
        RECT  2.840 4.640 3.960 5.440 ;
        RECT  3.960 3.990 3.970 5.440 ;
        RECT  3.970 3.790 4.370 5.440 ;
        RECT  4.370 3.990 4.380 5.440 ;
        RECT  4.380 4.640 5.510 5.440 ;
        RECT  5.510 3.990 5.520 5.440 ;
        RECT  5.520 3.790 5.920 5.440 ;
        RECT  5.920 3.990 5.930 5.440 ;
        RECT  5.930 4.640 7.050 5.440 ;
        RECT  7.050 4.310 7.060 5.440 ;
        RECT  7.060 4.110 7.460 5.440 ;
        RECT  7.460 4.310 7.470 5.440 ;
        RECT  7.470 4.640 8.640 5.440 ;
        RECT  8.640 3.260 8.650 5.440 ;
        RECT  8.650 3.060 9.050 5.440 ;
        RECT  9.050 3.260 9.060 5.440 ;
        RECT  9.060 4.640 9.240 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.240 0.400 ;
        RECT  1.240 -0.400 1.250 0.850 ;
        RECT  1.250 -0.400 1.650 1.050 ;
        RECT  1.650 -0.400 1.660 0.850 ;
        RECT  1.660 -0.400 2.660 0.400 ;
        RECT  2.660 -0.400 3.060 0.930 ;
        RECT  3.060 -0.400 4.030 0.400 ;
        RECT  4.030 -0.400 4.040 0.730 ;
        RECT  4.040 -0.400 4.440 0.930 ;
        RECT  4.440 -0.400 4.450 0.730 ;
        RECT  4.450 -0.400 5.530 0.400 ;
        RECT  5.530 -0.400 5.540 0.730 ;
        RECT  5.540 -0.400 5.940 0.930 ;
        RECT  5.940 -0.400 5.950 0.730 ;
        RECT  5.950 -0.400 7.000 0.400 ;
        RECT  7.000 -0.400 7.010 0.730 ;
        RECT  7.010 -0.400 7.410 0.930 ;
        RECT  7.410 -0.400 7.420 0.730 ;
        RECT  7.420 -0.400 9.240 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.910 2.160 6.470 2.560 ;
        RECT  2.930 2.150 4.910 2.570 ;
        RECT  2.510 1.380 2.930 3.340 ;
        RECT  0.830 1.380 2.510 1.800 ;
        RECT  0.370 2.920 2.510 3.340 ;
        RECT  0.630 1.390 0.830 1.790 ;
        RECT  0.170 2.930 0.370 3.330 ;
    END
END BUFX16

MACRO BUFX12
    CLASS CORE ;
    FOREIGN BUFX12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ BUFXL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.860 2.830 4.830 3.510 ;
        RECT  2.750 1.140 4.830 1.820 ;
        RECT  4.830 1.140 6.390 3.510 ;
        RECT  6.390 1.140 6.400 1.390 ;
        RECT  6.390 2.510 6.490 3.510 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.660 1.840 0.860 2.370 ;
        RECT  0.860 1.830 1.120 2.370 ;
        RECT  1.120 1.960 1.130 2.370 ;
        RECT  1.130 1.960 1.210 2.360 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.780 5.440 ;
        RECT  0.780 3.850 0.790 5.440 ;
        RECT  0.790 3.650 1.190 5.440 ;
        RECT  1.190 3.850 1.200 5.440 ;
        RECT  1.200 4.640 2.240 5.440 ;
        RECT  2.240 4.210 2.250 5.440 ;
        RECT  2.250 4.010 2.650 5.440 ;
        RECT  2.650 4.210 2.660 5.440 ;
        RECT  2.660 4.640 3.760 5.440 ;
        RECT  3.760 4.210 3.770 5.440 ;
        RECT  3.770 4.010 4.170 5.440 ;
        RECT  4.170 4.210 4.180 5.440 ;
        RECT  4.180 4.640 5.300 5.440 ;
        RECT  5.300 4.210 5.310 5.440 ;
        RECT  5.310 4.010 5.710 5.440 ;
        RECT  5.710 4.210 5.720 5.440 ;
        RECT  5.720 4.640 6.690 5.440 ;
        RECT  6.690 4.210 6.700 5.440 ;
        RECT  6.700 4.010 7.100 5.440 ;
        RECT  7.100 4.210 7.110 5.440 ;
        RECT  7.110 4.640 7.920 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.820 0.400 ;
        RECT  0.820 -0.400 1.220 0.560 ;
        RECT  1.220 -0.400 2.240 0.400 ;
        RECT  2.240 -0.400 2.250 0.670 ;
        RECT  2.250 -0.400 2.650 0.870 ;
        RECT  2.650 -0.400 2.660 0.670 ;
        RECT  2.660 -0.400 3.550 0.400 ;
        RECT  3.550 -0.400 3.560 0.670 ;
        RECT  3.560 -0.400 3.960 0.870 ;
        RECT  3.960 -0.400 3.970 0.670 ;
        RECT  3.970 -0.400 4.890 0.400 ;
        RECT  4.890 -0.400 4.900 0.670 ;
        RECT  4.900 -0.400 5.300 0.870 ;
        RECT  5.300 -0.400 5.310 0.670 ;
        RECT  5.310 -0.400 6.180 0.400 ;
        RECT  6.180 -0.400 6.190 0.670 ;
        RECT  6.190 -0.400 6.590 0.870 ;
        RECT  6.590 -0.400 6.600 0.670 ;
        RECT  6.600 -0.400 7.920 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.730 2.150 4.500 2.550 ;
        RECT  1.900 2.140 3.730 2.560 ;
        RECT  1.890 1.590 1.900 3.160 ;
        RECT  1.490 1.390 1.890 3.160 ;
        RECT  1.480 1.590 1.490 3.160 ;
        RECT  0.370 2.740 1.480 3.160 ;
        RECT  0.170 2.750 0.370 3.150 ;
    END
END BUFX12

MACRO AOI33XL
    CLASS CORE ;
    FOREIGN AOI33XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.080 1.020 2.480 1.420 ;
        RECT  3.040 3.110 3.200 3.510 ;
        RECT  3.200 3.010 3.440 3.510 ;
        RECT  3.440 3.010 4.560 3.250 ;
        RECT  4.560 3.010 4.830 3.510 ;
        RECT  4.820 2.390 4.830 2.650 ;
        RECT  2.480 1.020 4.830 1.260 ;
        RECT  4.830 1.020 4.960 3.510 ;
        RECT  4.960 1.020 5.070 3.250 ;
        RECT  5.070 2.390 5.080 2.650 ;
        END
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.810 0.520 2.420 ;
        RECT  0.520 1.820 0.550 2.420 ;
        RECT  0.550 1.820 0.890 2.220 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 1.120 3.210 ;
        RECT  1.120 2.950 1.180 3.190 ;
        RECT  1.180 2.540 1.420 3.190 ;
        RECT  1.420 2.540 1.580 2.940 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.790 2.090 ;
        RECT  1.790 1.750 2.190 2.150 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.030 1.610 4.040 1.930 ;
        RECT  4.040 1.610 4.120 2.070 ;
        RECT  4.120 1.610 4.160 2.080 ;
        RECT  4.160 1.610 4.420 2.090 ;
        RECT  4.420 1.610 4.440 2.070 ;
        RECT  4.440 1.610 4.450 1.930 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.240 2.270 3.640 2.670 ;
        RECT  3.640 2.390 3.760 2.650 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 2.950 2.440 3.210 ;
        RECT  2.440 2.950 2.530 3.190 ;
        RECT  2.530 2.290 2.770 3.190 ;
        RECT  2.770 2.290 2.930 2.690 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.670 5.440 ;
        RECT  1.670 4.480 2.070 5.440 ;
        RECT  2.070 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.310 0.400 ;
        RECT  0.310 -0.400 0.710 0.560 ;
        RECT  0.710 -0.400 3.980 0.400 ;
        RECT  3.980 -0.400 4.380 0.560 ;
        RECT  4.380 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.040 3.490 4.200 3.890 ;
        RECT  3.800 3.490 4.040 3.990 ;
        RECT  2.690 3.750 3.800 3.990 ;
        RECT  2.670 3.490 2.690 3.990 ;
        RECT  2.290 3.490 2.670 4.030 ;
        RECT  1.240 3.790 2.290 4.030 ;
        RECT  0.840 3.570 1.240 4.030 ;
    END
END AOI33XL

MACRO AOI33X4
    CLASS CORE ;
    FOREIGN AOI33X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI33XL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.710 1.170 7.140 3.220 ;
        RECT  7.140 1.820 7.150 3.220 ;
        END
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.460 2.420 ;
        RECT  0.460 1.840 0.500 2.420 ;
        RECT  0.500 1.840 0.540 2.410 ;
        RECT  0.540 2.010 0.870 2.410 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 1.200 3.210 ;
        RECT  1.200 2.810 1.600 3.210 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.670 2.090 ;
        RECT  1.670 1.820 2.070 2.220 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.080 2.390 4.520 2.820 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.510 2.090 ;
        RECT  3.510 1.830 3.750 2.810 ;
        RECT  3.750 1.830 3.760 2.090 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.710 2.930 2.850 3.170 ;
        RECT  2.840 2.390 2.850 2.650 ;
        RECT  2.850 2.390 3.090 3.170 ;
        RECT  3.090 2.390 3.100 2.650 ;
        RECT  3.090 2.930 3.110 3.170 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.190 5.440 ;
        RECT  0.190 4.130 0.200 5.440 ;
        RECT  0.200 3.930 0.600 5.440 ;
        RECT  0.600 4.130 0.610 5.440 ;
        RECT  0.610 4.640 1.700 5.440 ;
        RECT  1.700 4.010 2.100 5.440 ;
        RECT  2.100 4.640 6.090 5.440 ;
        RECT  6.090 4.010 6.490 5.440 ;
        RECT  6.490 4.640 7.360 5.440 ;
        RECT  7.360 4.010 7.760 5.440 ;
        RECT  7.760 4.640 7.920 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 3.640 0.400 ;
        RECT  3.640 -0.400 3.650 0.900 ;
        RECT  3.650 -0.400 4.050 1.020 ;
        RECT  4.050 -0.400 4.060 0.900 ;
        RECT  4.060 -0.400 6.030 0.400 ;
        RECT  6.030 -0.400 6.040 0.690 ;
        RECT  6.040 -0.400 6.440 0.890 ;
        RECT  6.440 -0.400 6.450 0.690 ;
        RECT  6.450 -0.400 7.340 0.400 ;
        RECT  7.340 -0.400 7.350 0.690 ;
        RECT  7.350 -0.400 7.750 0.890 ;
        RECT  7.750 -0.400 7.760 0.690 ;
        RECT  7.760 -0.400 7.920 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.200 1.310 6.440 3.250 ;
        RECT  5.650 1.310 6.200 1.550 ;
        RECT  5.570 3.010 6.200 3.250 ;
        RECT  5.030 1.930 5.800 2.170 ;
        RECT  5.410 0.670 5.650 1.550 ;
        RECT  5.330 3.010 5.570 3.410 ;
        RECT  5.250 0.670 5.410 0.910 ;
        RECT  5.030 3.830 5.050 4.070 ;
        RECT  4.790 1.300 5.030 4.070 ;
        RECT  2.310 1.300 4.790 1.540 ;
        RECT  4.650 3.220 4.790 4.070 ;
        RECT  4.640 3.220 4.650 3.860 ;
        RECT  3.630 3.220 4.640 3.460 ;
        RECT  3.930 3.750 4.330 4.360 ;
        RECT  2.880 4.120 3.930 4.360 ;
        RECT  3.390 3.220 3.630 3.770 ;
        RECT  3.210 3.530 3.390 3.770 ;
        RECT  2.730 3.490 2.880 4.360 ;
        RECT  2.470 3.490 2.730 4.370 ;
        RECT  1.340 3.490 2.470 3.730 ;
        RECT  2.460 4.090 2.470 4.370 ;
        RECT  1.910 1.100 2.310 1.540 ;
        RECT  0.940 3.490 1.340 4.090 ;
    END
END AOI33X4

MACRO AOI33X2
    CLASS CORE ;
    FOREIGN AOI33X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI33XL ;
    SIZE 9.240 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.900 0.730 3.090 0.970 ;
        RECT  3.090 0.730 3.330 1.340 ;
        RECT  3.330 1.100 5.390 1.340 ;
        RECT  5.390 0.960 5.550 1.340 ;
        RECT  5.550 0.800 5.950 1.340 ;
        RECT  4.870 3.040 7.950 3.440 ;
        RECT  7.950 3.040 8.790 3.280 ;
        RECT  8.780 2.390 8.790 2.650 ;
        RECT  5.950 1.100 8.790 1.340 ;
        RECT  8.790 1.100 9.030 3.280 ;
        RECT  9.030 2.390 9.040 2.650 ;
        END
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.410 2.650 ;
        RECT  0.410 2.390 0.460 2.990 ;
        RECT  0.460 2.400 0.650 2.990 ;
        RECT  0.650 2.590 0.810 2.990 ;
        RECT  0.810 2.670 3.410 2.910 ;
        RECT  3.410 2.270 3.810 2.910 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 1.120 2.090 ;
        RECT  1.120 1.850 1.130 2.090 ;
        RECT  1.130 1.850 1.370 2.380 ;
        RECT  1.370 1.970 1.530 2.380 ;
        RECT  1.530 2.140 2.600 2.380 ;
        RECT  2.600 1.970 3.000 2.380 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.880 1.390 2.090 1.860 ;
        RECT  2.090 1.290 2.180 1.860 ;
        RECT  2.180 1.270 2.330 1.860 ;
        RECT  2.330 1.270 2.440 1.530 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.130 1.620 4.160 2.020 ;
        RECT  4.160 1.620 4.420 2.090 ;
        RECT  4.420 1.620 4.530 2.020 ;
        RECT  4.530 1.700 7.680 1.940 ;
        RECT  7.680 1.620 8.080 2.020 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.820 2.280 5.450 2.660 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.850 2.380 5.860 2.660 ;
        RECT  5.860 2.220 6.260 2.660 ;
        RECT  6.260 2.380 6.570 2.660 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.770 5.440 ;
        RECT  0.770 4.150 0.780 5.440 ;
        RECT  0.780 3.950 1.180 5.440 ;
        RECT  1.180 4.150 1.190 5.440 ;
        RECT  1.190 4.640 2.120 5.440 ;
        RECT  2.120 4.150 2.130 5.440 ;
        RECT  2.130 3.950 2.530 5.440 ;
        RECT  2.530 4.150 2.540 5.440 ;
        RECT  2.540 4.640 3.460 5.440 ;
        RECT  3.460 4.150 3.470 5.440 ;
        RECT  3.470 3.950 3.870 5.440 ;
        RECT  3.870 4.150 3.880 5.440 ;
        RECT  3.880 4.640 9.240 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.230 0.400 ;
        RECT  0.230 -0.400 0.240 0.790 ;
        RECT  0.240 -0.400 0.640 0.990 ;
        RECT  0.640 -0.400 0.650 0.790 ;
        RECT  0.650 -0.400 3.730 0.400 ;
        RECT  3.730 -0.400 4.130 0.560 ;
        RECT  4.130 -0.400 7.300 0.400 ;
        RECT  7.300 -0.400 7.700 0.560 ;
        RECT  7.700 -0.400 9.240 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  8.370 3.720 8.570 4.120 ;
        RECT  4.560 3.710 8.370 4.130 ;
        RECT  4.140 3.260 4.560 4.130 ;
        RECT  0.370 3.260 4.140 3.680 ;
        RECT  0.170 3.270 0.370 3.670 ;
    END
END AOI33X2

MACRO AOI33X1
    CLASS CORE ;
    FOREIGN AOI33X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI33XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.080 0.820 2.480 1.220 ;
        RECT  3.040 3.060 3.440 3.490 ;
        RECT  3.440 3.060 4.560 3.300 ;
        RECT  2.480 0.980 4.730 1.220 ;
        RECT  4.560 3.060 4.810 3.490 ;
        RECT  4.810 3.060 4.830 3.500 ;
        RECT  4.820 2.390 4.830 2.650 ;
        RECT  4.730 0.980 4.830 1.260 ;
        RECT  4.830 0.980 5.070 3.500 ;
        RECT  5.070 3.200 5.080 3.500 ;
        RECT  5.070 2.390 5.080 2.650 ;
        END
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.550 2.420 ;
        RECT  0.550 1.830 0.640 2.250 ;
        RECT  0.640 1.830 1.010 2.240 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 1.190 3.210 ;
        RECT  1.190 2.860 1.590 3.260 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.630 2.090 ;
        RECT  1.630 1.820 1.790 2.090 ;
        RECT  1.790 1.820 2.190 2.220 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.050 1.610 4.160 2.010 ;
        RECT  4.160 1.610 4.420 2.090 ;
        RECT  4.420 1.610 4.450 2.010 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.240 2.270 3.640 2.670 ;
        RECT  3.640 2.390 3.760 2.650 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 2.950 2.440 3.210 ;
        RECT  2.440 2.950 2.530 3.190 ;
        RECT  2.530 2.260 2.770 3.190 ;
        RECT  2.770 2.260 2.930 2.660 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.190 0.180 5.440 ;
        RECT  0.180 3.990 0.580 5.440 ;
        RECT  0.580 4.190 0.590 5.440 ;
        RECT  0.590 4.640 1.760 5.440 ;
        RECT  1.760 4.480 2.160 5.440 ;
        RECT  2.160 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.310 0.400 ;
        RECT  0.310 -0.400 0.710 0.560 ;
        RECT  0.710 -0.400 3.980 0.400 ;
        RECT  3.980 -0.400 4.380 0.560 ;
        RECT  4.380 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.800 3.580 4.200 4.010 ;
        RECT  2.680 3.770 3.800 4.010 ;
        RECT  2.280 3.580 2.680 4.010 ;
        RECT  1.340 3.770 2.280 4.010 ;
        RECT  0.940 3.580 1.340 4.010 ;
    END
END AOI33X1

MACRO AOI32XL
    CLASS CORE ;
    FOREIGN AOI32XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.900 1.160 1.910 1.550 ;
        RECT  1.910 0.800 2.180 1.550 ;
        RECT  2.180 0.800 2.310 1.540 ;
        RECT  3.220 2.940 3.230 3.420 ;
        RECT  3.230 2.940 3.620 3.560 ;
        RECT  3.620 2.950 3.630 3.560 ;
        RECT  3.630 2.950 4.170 3.190 ;
        RECT  4.160 2.390 4.170 2.650 ;
        RECT  2.310 1.300 4.170 1.540 ;
        RECT  4.170 1.300 4.410 3.190 ;
        RECT  4.410 2.390 4.420 2.650 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.760 2.420 ;
        RECT  3.760 1.840 3.800 2.420 ;
        RECT  3.800 2.040 3.810 2.420 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.730 2.180 2.840 2.580 ;
        RECT  2.840 2.180 3.100 2.650 ;
        RECT  3.100 2.180 3.130 2.640 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.460 2.420 ;
        RECT  0.460 1.840 0.500 2.420 ;
        RECT  0.500 1.840 0.540 2.410 ;
        RECT  0.540 2.010 0.870 2.410 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 1.120 3.210 ;
        RECT  1.120 2.950 1.200 3.190 ;
        RECT  1.200 2.540 1.440 3.190 ;
        RECT  1.440 2.540 1.600 3.090 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.680 2.090 ;
        RECT  1.680 1.820 2.080 2.220 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.190 0.180 5.440 ;
        RECT  0.180 3.990 0.580 5.440 ;
        RECT  0.580 4.190 0.590 5.440 ;
        RECT  0.590 4.640 1.700 5.440 ;
        RECT  1.700 4.070 2.100 5.440 ;
        RECT  2.100 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 3.190 0.400 ;
        RECT  3.190 -0.400 3.590 0.560 ;
        RECT  3.590 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.990 3.610 4.390 4.080 ;
        RECT  2.880 3.840 3.990 4.080 ;
        RECT  2.470 3.550 2.880 4.080 ;
        RECT  1.340 3.550 2.470 3.790 ;
        RECT  0.940 3.550 1.340 4.010 ;
    END
END AOI32XL

MACRO AOI32X4
    CLASS CORE ;
    FOREIGN AOI32X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI32XL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  5.970 2.750 6.050 3.150 ;
        RECT  5.920 1.270 6.050 1.670 ;
        RECT  6.050 1.270 6.320 3.220 ;
        RECT  6.320 1.820 6.490 3.220 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.890 1.820 3.500 2.060 ;
        RECT  3.500 1.820 3.750 2.090 ;
        RECT  3.750 1.830 3.760 2.090 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.640 2.390 3.120 2.870 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.460 2.420 ;
        RECT  0.460 1.840 0.500 2.420 ;
        RECT  0.500 1.840 0.540 2.410 ;
        RECT  0.540 2.010 0.870 2.410 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 1.200 3.210 ;
        RECT  1.200 2.810 1.600 3.210 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.680 2.090 ;
        RECT  1.680 1.820 2.080 2.220 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.130 0.180 5.440 ;
        RECT  0.180 3.930 0.580 5.440 ;
        RECT  0.580 4.130 0.590 5.440 ;
        RECT  0.590 4.640 1.700 5.440 ;
        RECT  1.700 4.010 2.100 5.440 ;
        RECT  2.100 4.640 5.310 5.440 ;
        RECT  5.310 4.010 5.710 5.440 ;
        RECT  5.710 4.640 6.620 5.440 ;
        RECT  6.620 4.010 7.020 5.440 ;
        RECT  7.020 4.640 7.260 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 3.180 0.400 ;
        RECT  3.180 -0.400 3.190 0.900 ;
        RECT  3.190 -0.400 3.590 1.020 ;
        RECT  3.590 -0.400 3.600 0.900 ;
        RECT  3.600 -0.400 5.240 0.400 ;
        RECT  5.240 -0.400 5.250 0.790 ;
        RECT  5.250 -0.400 5.650 0.990 ;
        RECT  5.650 -0.400 5.660 0.790 ;
        RECT  5.660 -0.400 6.560 0.400 ;
        RECT  6.560 -0.400 6.570 0.790 ;
        RECT  6.570 -0.400 6.970 0.990 ;
        RECT  6.970 -0.400 6.980 0.790 ;
        RECT  6.980 -0.400 7.260 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.580 2.030 5.770 2.430 ;
        RECT  5.340 1.410 5.580 3.330 ;
        RECT  4.890 1.410 5.340 1.650 ;
        RECT  4.490 3.090 5.340 3.330 ;
        RECT  4.360 1.930 5.060 2.170 ;
        RECT  4.650 0.720 4.890 1.650 ;
        RECT  4.490 0.720 4.650 0.960 ;
        RECT  3.990 3.750 4.390 4.360 ;
        RECT  4.120 1.300 4.360 2.620 ;
        RECT  2.310 1.300 4.120 1.540 ;
        RECT  3.710 2.380 4.120 2.620 ;
        RECT  2.880 4.120 3.990 4.360 ;
        RECT  3.470 2.380 3.710 3.770 ;
        RECT  3.230 3.530 3.470 3.770 ;
        RECT  2.730 3.490 2.880 4.360 ;
        RECT  2.470 3.490 2.730 4.370 ;
        RECT  1.340 3.490 2.470 3.730 ;
        RECT  2.460 4.090 2.470 4.370 ;
        RECT  1.910 1.100 2.310 1.540 ;
        RECT  0.940 3.490 1.340 4.090 ;
    END
END AOI32X4

MACRO AOI32X2
    CLASS CORE ;
    FOREIGN AOI32X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI32XL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.570 0.750 3.230 0.990 ;
        RECT  3.230 0.750 3.470 1.550 ;
        RECT  3.470 1.280 3.510 1.550 ;
        RECT  3.510 1.310 5.590 1.550 ;
        RECT  5.590 0.860 6.150 1.550 ;
        RECT  5.330 3.100 6.990 3.500 ;
        RECT  6.990 3.100 7.470 3.340 ;
        RECT  7.460 2.390 7.470 2.650 ;
        RECT  6.150 1.310 7.470 1.550 ;
        RECT  7.470 1.310 7.710 3.340 ;
        RECT  7.710 2.390 7.720 2.650 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.790 1.850 4.820 2.090 ;
        RECT  4.820 1.830 4.950 2.090 ;
        RECT  4.950 1.830 5.080 2.760 ;
        RECT  5.080 1.850 5.190 2.760 ;
        RECT  5.190 2.520 6.670 2.760 ;
        RECT  6.670 2.420 7.070 2.820 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.830 1.800 6.430 2.200 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 0.890 2.650 ;
        RECT  0.890 2.390 1.120 2.910 ;
        RECT  1.120 2.410 1.210 2.910 ;
        RECT  1.210 2.670 4.180 2.910 ;
        RECT  4.180 2.610 4.580 2.910 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.660 1.970 1.900 2.380 ;
        RECT  1.900 2.140 3.270 2.380 ;
        RECT  3.270 1.840 3.500 2.380 ;
        RECT  3.500 1.830 3.670 2.380 ;
        RECT  3.670 1.830 3.760 2.090 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 1.270 2.290 1.530 ;
        RECT  2.290 1.270 2.440 1.860 ;
        RECT  2.440 1.290 2.530 1.860 ;
        RECT  2.530 1.620 2.950 1.860 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.170 5.440 ;
        RECT  1.170 4.150 1.180 5.440 ;
        RECT  1.180 3.950 1.580 5.440 ;
        RECT  1.580 4.150 1.590 5.440 ;
        RECT  1.590 4.640 2.510 5.440 ;
        RECT  2.510 4.150 2.520 5.440 ;
        RECT  2.520 3.950 2.920 5.440 ;
        RECT  2.920 4.150 2.930 5.440 ;
        RECT  2.930 4.640 3.850 5.440 ;
        RECT  3.850 4.150 3.860 5.440 ;
        RECT  3.860 3.950 4.260 5.440 ;
        RECT  4.260 4.150 4.270 5.440 ;
        RECT  4.270 4.640 7.920 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.900 0.400 ;
        RECT  0.900 -0.400 0.910 0.790 ;
        RECT  0.910 -0.400 1.310 0.990 ;
        RECT  1.310 -0.400 1.320 0.790 ;
        RECT  1.320 -0.400 4.300 0.400 ;
        RECT  4.300 -0.400 4.310 0.830 ;
        RECT  4.310 -0.400 4.710 1.030 ;
        RECT  4.710 -0.400 4.720 0.830 ;
        RECT  4.720 -0.400 6.970 0.400 ;
        RECT  6.970 -0.400 6.980 0.830 ;
        RECT  6.980 -0.400 7.380 0.950 ;
        RECT  7.380 -0.400 7.390 0.830 ;
        RECT  7.390 -0.400 7.920 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  7.430 3.780 7.630 4.180 ;
        RECT  5.040 3.770 7.430 4.190 ;
        RECT  4.830 3.260 5.040 4.190 ;
        RECT  4.630 3.260 4.830 4.180 ;
        RECT  4.620 3.260 4.630 3.980 ;
        RECT  0.760 3.260 4.620 3.680 ;
        RECT  0.560 3.270 0.760 3.670 ;
    END
END AOI32X2

MACRO AOI32X1
    CLASS CORE ;
    FOREIGN AOI32X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI32XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.910 1.040 2.310 1.540 ;
        RECT  3.230 3.090 3.630 3.490 ;
        RECT  3.630 3.090 4.170 3.330 ;
        RECT  4.160 2.390 4.170 2.650 ;
        RECT  2.310 1.300 4.170 1.540 ;
        RECT  4.170 1.300 4.410 3.330 ;
        RECT  4.410 2.390 4.420 2.650 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.760 2.420 ;
        RECT  3.760 1.840 3.800 2.420 ;
        RECT  3.800 2.040 3.810 2.420 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.730 2.180 2.840 2.580 ;
        RECT  2.840 2.180 3.100 2.650 ;
        RECT  3.100 2.180 3.130 2.640 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.460 2.420 ;
        RECT  0.460 1.840 0.520 2.420 ;
        RECT  0.520 1.840 0.540 2.410 ;
        RECT  0.540 2.010 0.890 2.410 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 1.120 3.210 ;
        RECT  1.120 2.950 1.210 3.190 ;
        RECT  1.210 2.540 1.480 3.190 ;
        RECT  1.480 2.540 1.640 3.080 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.680 2.090 ;
        RECT  1.680 1.820 2.080 2.220 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.190 0.180 5.440 ;
        RECT  0.180 3.990 0.580 5.440 ;
        RECT  0.580 4.190 0.590 5.440 ;
        RECT  0.590 4.640 1.690 5.440 ;
        RECT  1.690 4.130 1.700 5.440 ;
        RECT  1.700 4.010 2.100 5.440 ;
        RECT  2.100 4.130 2.110 5.440 ;
        RECT  2.110 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 3.120 0.400 ;
        RECT  3.120 -0.400 3.130 0.900 ;
        RECT  3.130 -0.400 3.530 1.020 ;
        RECT  3.530 -0.400 3.540 0.900 ;
        RECT  3.540 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.990 3.730 4.390 4.150 ;
        RECT  2.880 3.910 3.990 4.150 ;
        RECT  2.640 3.490 2.880 4.150 ;
        RECT  2.470 3.490 2.640 3.910 ;
        RECT  1.340 3.490 2.470 3.730 ;
        RECT  0.940 3.490 1.340 3.910 ;
    END
END AOI32X1

MACRO AOI31XL
    CLASS CORE ;
    FOREIGN AOI31XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.910 1.090 2.310 1.490 ;
        RECT  3.330 2.970 3.510 3.370 ;
        RECT  3.500 2.390 3.510 2.650 ;
        RECT  2.310 1.250 3.510 1.490 ;
        RECT  3.510 1.250 3.750 3.370 ;
        RECT  3.750 2.390 3.760 2.650 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 1.830 2.900 2.090 ;
        RECT  2.900 1.830 3.100 2.580 ;
        RECT  3.100 1.850 3.140 2.580 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.220 2.090 ;
        RECT  0.220 1.830 0.410 2.580 ;
        RECT  0.410 1.830 0.460 2.740 ;
        RECT  0.460 2.340 0.810 2.740 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 1.050 2.090 ;
        RECT  1.050 1.830 1.120 2.640 ;
        RECT  1.120 1.840 1.290 2.640 ;
        RECT  1.290 2.400 1.530 2.640 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.890 1.870 2.050 2.270 ;
        RECT  2.050 1.870 2.180 2.630 ;
        RECT  2.180 1.870 2.290 2.650 ;
        RECT  2.290 2.390 2.440 2.650 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 3.350 0.570 5.440 ;
        RECT  0.570 4.640 1.740 5.440 ;
        RECT  1.740 3.690 1.750 5.440 ;
        RECT  1.750 3.570 2.150 5.440 ;
        RECT  2.150 3.690 2.160 5.440 ;
        RECT  2.160 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 2.780 0.400 ;
        RECT  2.780 -0.400 2.790 0.770 ;
        RECT  2.790 -0.400 3.190 0.890 ;
        RECT  3.190 -0.400 3.200 0.770 ;
        RECT  3.200 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.570 2.970 2.970 3.370 ;
        RECT  1.330 3.060 2.570 3.300 ;
        RECT  0.930 2.980 1.330 3.380 ;
    END
END AOI31XL

MACRO AOI31X4
    CLASS CORE ;
    FOREIGN AOI31X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI31XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.920 2.880 5.320 3.840 ;
        RECT  5.320 2.880 5.390 3.780 ;
        RECT  5.390 2.380 5.580 3.780 ;
        RECT  4.850 1.220 5.580 1.460 ;
        RECT  5.580 1.220 5.820 3.780 ;
        RECT  5.820 2.380 5.830 3.780 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.750 1.560 3.200 2.100 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.860 0.510 2.650 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 1.380 3.010 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 1.820 1.680 2.100 ;
        RECT  1.680 1.820 1.920 2.350 ;
        RECT  1.920 1.820 1.930 2.100 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.380 5.440 ;
        RECT  1.380 4.480 1.780 5.440 ;
        RECT  1.780 4.640 4.140 5.440 ;
        RECT  4.140 4.250 4.150 5.440 ;
        RECT  4.150 4.050 4.550 5.440 ;
        RECT  4.550 4.250 4.560 5.440 ;
        RECT  4.560 4.640 5.560 5.440 ;
        RECT  5.560 4.370 5.570 5.440 ;
        RECT  5.570 4.170 5.970 5.440 ;
        RECT  5.970 4.370 5.980 5.440 ;
        RECT  5.980 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 1.260 ;
        RECT  0.570 -0.400 2.720 0.400 ;
        RECT  2.720 -0.400 2.730 1.090 ;
        RECT  2.730 -0.400 3.130 1.290 ;
        RECT  3.130 -0.400 3.140 1.090 ;
        RECT  3.140 -0.400 4.200 0.400 ;
        RECT  4.200 -0.400 4.210 0.700 ;
        RECT  4.210 -0.400 4.610 0.900 ;
        RECT  4.610 -0.400 4.620 0.700 ;
        RECT  4.620 -0.400 5.480 0.400 ;
        RECT  5.480 -0.400 5.490 0.700 ;
        RECT  5.490 -0.400 5.890 0.900 ;
        RECT  5.890 -0.400 5.900 0.700 ;
        RECT  5.900 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.790 1.780 5.120 2.180 ;
        RECT  4.520 1.770 4.790 2.190 ;
        RECT  4.280 1.180 4.520 3.680 ;
        RECT  3.870 1.180 4.280 1.420 ;
        RECT  3.830 3.440 4.280 3.680 ;
        RECT  3.600 2.220 4.000 2.620 ;
        RECT  3.630 1.000 3.870 1.420 ;
        RECT  3.430 3.440 3.830 3.840 ;
        RECT  3.470 1.000 3.630 1.400 ;
        RECT  3.310 2.380 3.600 2.620 ;
        RECT  2.910 2.380 3.310 3.100 ;
        RECT  2.900 2.380 2.910 2.740 ;
        RECT  2.450 2.380 2.900 2.620 ;
        RECT  2.410 3.000 2.570 3.400 ;
        RECT  2.250 1.110 2.450 2.620 ;
        RECT  2.170 3.000 2.410 3.730 ;
        RECT  2.210 0.950 2.250 2.620 ;
        RECT  1.850 0.950 2.210 1.350 ;
        RECT  1.170 3.490 2.170 3.730 ;
        RECT  0.770 3.490 1.170 3.890 ;
    END
END AOI31X4

MACRO AOI31X2
    CLASS CORE ;
    FOREIGN AOI31X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI31XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.330 0.750 1.480 0.990 ;
        RECT  1.480 0.750 1.720 1.390 ;
        RECT  1.720 0.960 1.770 1.390 ;
        RECT  1.770 1.150 3.750 1.390 ;
        RECT  3.750 1.150 3.900 1.540 ;
        RECT  3.900 0.660 4.180 1.620 ;
        RECT  4.180 0.660 4.300 2.900 ;
        RECT  4.300 1.270 4.420 2.900 ;
        RECT  4.420 2.660 4.730 2.900 ;
        RECT  4.730 2.660 4.860 2.960 ;
        RECT  4.860 2.660 5.100 3.500 ;
        RECT  5.100 3.100 5.260 3.500 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.820 1.830 4.830 2.090 ;
        RECT  4.830 1.830 5.080 2.380 ;
        RECT  5.080 1.980 5.260 2.380 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.270 0.970 1.530 ;
        RECT  0.970 1.270 1.120 1.910 ;
        RECT  1.120 1.290 1.210 1.910 ;
        RECT  1.210 1.670 2.470 1.910 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.190 2.190 2.750 2.430 ;
        RECT  2.750 2.050 2.840 2.430 ;
        RECT  2.840 1.830 2.990 2.430 ;
        RECT  2.990 1.830 3.100 2.370 ;
        RECT  3.100 1.970 3.280 2.370 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.460 2.650 ;
        RECT  0.460 2.410 0.550 2.650 ;
        RECT  0.550 2.410 0.560 2.660 ;
        RECT  0.560 2.410 0.800 2.950 ;
        RECT  0.800 2.710 3.680 2.950 ;
        RECT  3.680 2.100 3.920 2.950 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.780 5.440 ;
        RECT  0.780 3.980 0.790 5.440 ;
        RECT  0.790 3.780 1.190 5.440 ;
        RECT  1.190 3.980 1.200 5.440 ;
        RECT  1.200 4.640 2.120 5.440 ;
        RECT  2.120 3.980 2.130 5.440 ;
        RECT  2.130 3.780 2.530 5.440 ;
        RECT  2.530 3.980 2.540 5.440 ;
        RECT  2.540 4.640 3.460 5.440 ;
        RECT  3.460 3.980 3.470 5.440 ;
        RECT  3.470 3.780 3.870 5.440 ;
        RECT  3.870 3.980 3.880 5.440 ;
        RECT  3.880 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 2.090 0.400 ;
        RECT  2.090 -0.400 2.490 0.870 ;
        RECT  2.490 -0.400 4.770 0.400 ;
        RECT  4.770 -0.400 4.780 1.040 ;
        RECT  4.780 -0.400 5.180 1.520 ;
        RECT  5.180 -0.400 5.190 1.040 ;
        RECT  5.190 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.480 3.780 5.880 4.180 ;
        RECT  4.640 3.860 5.480 4.100 ;
        RECT  4.480 3.780 4.640 4.180 ;
        RECT  4.240 3.230 4.480 4.180 ;
        RECT  0.170 3.230 4.240 3.470 ;
    END
END AOI31X2

MACRO AOI31X1
    CLASS CORE ;
    FOREIGN AOI31X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI31XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.850 0.690 2.250 1.120 ;
        RECT  2.250 0.880 3.410 1.120 ;
        RECT  3.210 3.060 3.510 3.460 ;
        RECT  3.500 2.390 3.510 2.650 ;
        RECT  3.410 0.880 3.510 1.260 ;
        RECT  3.510 0.880 3.750 3.460 ;
        RECT  3.750 2.390 3.760 2.650 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.440 1.640 2.680 2.060 ;
        RECT  2.680 1.820 2.840 2.060 ;
        RECT  2.840 1.820 3.080 2.090 ;
        RECT  3.080 1.830 3.100 2.090 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.170 1.800 0.510 2.620 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 1.120 2.440 ;
        RECT  1.120 1.840 1.320 2.440 ;
        RECT  1.320 1.840 1.470 2.430 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.000 2.390 2.530 2.920 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.000 0.170 5.440 ;
        RECT  0.170 3.800 0.570 5.440 ;
        RECT  0.570 4.000 0.580 5.440 ;
        RECT  0.580 4.640 1.690 5.440 ;
        RECT  1.690 3.800 2.090 5.440 ;
        RECT  2.090 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 0.670 ;
        RECT  0.170 -0.400 0.570 0.790 ;
        RECT  0.570 -0.400 0.580 0.670 ;
        RECT  0.580 -0.400 2.670 0.400 ;
        RECT  2.670 -0.400 3.070 0.560 ;
        RECT  3.070 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  0.930 3.280 2.850 3.520 ;
    END
END AOI31X1

MACRO AOI2BB2XL
    CLASS CORE ;
    FOREIGN AOI2BB2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 2.950 3.510 3.210 ;
        RECT  2.990 1.380 3.510 1.620 ;
        RECT  3.510 1.380 3.750 3.210 ;
        RECT  3.750 2.950 3.760 3.210 ;
        RECT  3.760 2.960 3.770 3.210 ;
        RECT  3.770 2.960 4.010 4.130 ;
        RECT  4.010 3.730 4.170 4.130 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.000 1.820 2.330 2.450 ;
        RECT  2.330 1.830 2.440 2.090 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.750 2.390 3.130 3.150 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.210 2.090 ;
        RECT  0.210 1.350 0.550 2.090 ;
        RECT  0.550 1.350 0.750 1.590 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.980 1.190 2.660 ;
        END
    END A0N
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 2.250 5.440 ;
        RECT  2.250 4.190 2.650 5.440 ;
        RECT  2.650 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 0.900 ;
        RECT  0.170 -0.400 0.570 1.020 ;
        RECT  0.570 -0.400 0.580 0.900 ;
        RECT  0.580 -0.400 1.920 0.400 ;
        RECT  1.920 -0.400 2.320 0.560 ;
        RECT  2.320 -0.400 3.860 0.400 ;
        RECT  3.860 -0.400 4.260 0.560 ;
        RECT  4.260 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.030 0.850 4.270 2.410 ;
        RECT  1.720 0.850 4.030 1.090 ;
        RECT  3.010 3.670 3.410 4.130 ;
        RECT  1.890 3.670 3.010 3.910 ;
        RECT  1.490 3.670 1.890 4.230 ;
        RECT  1.480 0.850 1.720 3.310 ;
        RECT  1.130 0.850 1.480 1.260 ;
        RECT  1.230 3.070 1.480 3.310 ;
    END
END AOI2BB2XL

MACRO AOI2BB2X4
    CLASS CORE ;
    FOREIGN AOI2BB2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI2BB2XL ;
    SIZE 10.560 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.030 3.970 3.150 4.370 ;
        RECT  3.150 2.760 3.230 4.370 ;
        RECT  3.230 2.760 3.390 4.380 ;
        RECT  3.430 0.660 3.670 1.620 ;
        RECT  3.670 0.830 3.850 1.620 ;
        RECT  3.390 2.760 4.070 3.000 ;
        RECT  3.850 1.200 4.070 1.620 ;
        RECT  4.070 2.500 4.100 3.000 ;
        RECT  4.070 1.200 4.100 1.960 ;
        RECT  4.100 1.200 4.340 3.000 ;
        RECT  3.390 3.960 4.650 4.380 ;
        RECT  4.650 3.970 4.850 4.370 ;
        RECT  4.340 1.200 5.350 1.440 ;
        RECT  5.350 0.770 5.750 1.440 ;
        RECT  5.750 0.840 5.830 1.440 ;
        RECT  5.830 1.200 7.710 1.440 ;
        RECT  7.710 0.970 7.720 1.450 ;
        RECT  7.720 0.770 8.120 1.450 ;
        RECT  8.120 0.970 8.130 1.450 ;
        RECT  8.130 1.030 8.690 1.450 ;
        RECT  8.690 0.700 9.130 2.100 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.820 1.830 4.830 2.090 ;
        RECT  4.830 1.720 5.160 2.090 ;
        RECT  5.160 1.720 5.560 2.470 ;
        RECT  5.560 1.720 7.590 1.960 ;
        RECT  7.590 1.720 7.900 2.100 ;
        RECT  7.900 1.720 8.140 2.640 ;
        RECT  8.140 2.400 9.130 2.640 ;
        RECT  9.130 2.400 9.530 2.800 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.140 2.390 6.230 2.650 ;
        RECT  6.230 2.360 7.630 2.760 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.260 2.330 0.500 3.740 ;
        RECT  0.500 3.500 2.000 3.740 ;
        RECT  2.000 1.900 2.240 3.740 ;
        RECT  2.240 2.950 2.440 3.210 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.770 1.720 1.210 2.200 ;
        END
    END A0N
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 2.300 5.440 ;
        RECT  2.300 4.480 2.700 5.440 ;
        RECT  2.700 4.640 6.000 5.440 ;
        RECT  6.000 3.960 6.010 5.440 ;
        RECT  6.010 3.760 6.410 5.440 ;
        RECT  6.410 3.960 6.420 5.440 ;
        RECT  6.420 4.640 7.560 5.440 ;
        RECT  7.560 3.960 7.570 5.440 ;
        RECT  7.570 3.760 7.970 5.440 ;
        RECT  7.970 3.960 7.980 5.440 ;
        RECT  7.980 4.640 9.120 5.440 ;
        RECT  9.120 3.960 9.130 5.440 ;
        RECT  9.130 3.760 9.530 5.440 ;
        RECT  9.530 3.960 9.540 5.440 ;
        RECT  9.540 4.640 10.560 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.790 0.400 ;
        RECT  0.790 -0.400 0.800 0.980 ;
        RECT  0.800 -0.400 1.200 1.460 ;
        RECT  1.200 -0.400 1.210 0.980 ;
        RECT  1.210 -0.400 2.520 0.400 ;
        RECT  2.520 -0.400 2.530 0.980 ;
        RECT  2.530 -0.400 2.930 1.100 ;
        RECT  2.930 -0.400 2.940 0.980 ;
        RECT  2.940 -0.400 4.110 0.400 ;
        RECT  4.110 -0.400 4.120 0.720 ;
        RECT  4.120 -0.400 4.520 0.920 ;
        RECT  4.520 -0.400 4.530 0.720 ;
        RECT  4.530 -0.400 6.530 0.400 ;
        RECT  6.530 -0.400 6.540 0.720 ;
        RECT  6.540 -0.400 6.940 0.920 ;
        RECT  6.940 -0.400 6.950 0.720 ;
        RECT  6.950 -0.400 10.560 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  10.050 3.080 10.250 3.480 ;
        RECT  5.620 3.070 10.050 3.490 ;
        RECT  5.570 3.070 5.620 3.680 ;
        RECT  5.150 3.070 5.570 3.690 ;
        RECT  3.870 3.270 5.150 3.690 ;
        RECT  3.670 3.280 3.870 3.680 ;
        RECT  3.420 1.890 3.820 2.290 ;
        RECT  2.760 1.890 3.420 2.130 ;
        RECT  2.520 1.380 2.760 2.130 ;
        RECT  2.110 1.380 2.520 1.620 ;
        RECT  1.720 0.780 2.110 1.620 ;
        RECT  1.710 0.780 1.720 3.220 ;
        RECT  1.480 1.380 1.710 3.220 ;
        RECT  1.230 2.980 1.480 3.220 ;
    END
END AOI2BB2X4

MACRO AOI2BB2X2
    CLASS CORE ;
    FOREIGN AOI2BB2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI2BB2XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.890 0.700 3.290 1.100 ;
        RECT  4.100 4.130 4.180 4.370 ;
        RECT  4.180 3.940 4.500 4.370 ;
        RECT  4.500 3.940 4.730 4.340 ;
        RECT  4.730 3.940 4.830 4.320 ;
        RECT  3.290 0.860 5.040 1.100 ;
        RECT  5.040 0.780 5.390 1.180 ;
        RECT  5.390 0.780 5.440 1.510 ;
        RECT  5.440 0.940 5.480 1.510 ;
        RECT  4.830 3.940 5.490 4.180 ;
        RECT  5.480 0.940 5.490 1.530 ;
        RECT  5.490 0.940 5.630 4.180 ;
        RECT  5.630 1.270 5.730 4.180 ;
        RECT  5.730 1.270 5.740 1.530 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.150 2.880 4.070 3.120 ;
        RECT  4.070 2.530 4.160 3.120 ;
        RECT  4.160 2.390 4.310 3.120 ;
        RECT  4.310 2.390 4.340 2.770 ;
        RECT  4.340 2.370 4.740 2.770 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.660 1.840 2.820 2.080 ;
        RECT  2.820 1.380 3.060 2.080 ;
        RECT  3.060 1.380 3.190 1.840 ;
        RECT  3.190 1.380 4.440 1.620 ;
        RECT  4.440 1.380 4.660 2.080 ;
        RECT  4.660 1.380 4.680 2.090 ;
        RECT  4.680 1.640 5.130 2.090 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.360 2.360 1.780 2.780 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.870 0.550 2.650 ;
        END
    END A0N
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.440 5.440 ;
        RECT  1.440 4.250 1.450 5.440 ;
        RECT  1.450 4.050 1.850 5.440 ;
        RECT  1.850 4.250 1.860 5.440 ;
        RECT  1.860 4.640 2.750 5.440 ;
        RECT  2.750 4.250 2.760 5.440 ;
        RECT  2.760 4.050 3.160 5.440 ;
        RECT  3.160 4.250 3.170 5.440 ;
        RECT  3.170 4.640 5.530 5.440 ;
        RECT  5.530 4.480 5.930 5.440 ;
        RECT  5.930 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.560 ;
        RECT  0.570 -0.400 1.420 0.400 ;
        RECT  1.420 -0.400 1.610 0.410 ;
        RECT  1.610 -0.400 2.010 1.460 ;
        RECT  2.010 -0.400 3.760 0.400 ;
        RECT  3.760 -0.400 4.160 0.560 ;
        RECT  4.160 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.830 3.400 5.200 3.640 ;
        RECT  3.510 3.400 3.830 3.690 ;
        RECT  3.460 1.900 3.700 2.600 ;
        RECT  2.090 3.450 3.510 3.690 ;
        RECT  2.380 2.360 3.460 2.600 ;
        RECT  2.140 1.810 2.380 2.600 ;
        RECT  1.250 1.810 2.140 2.050 ;
        RECT  1.060 1.180 1.250 2.050 ;
        RECT  0.820 1.180 1.060 3.320 ;
        RECT  0.570 3.080 0.820 3.320 ;
        RECT  0.170 3.080 0.570 3.480 ;
    END
END AOI2BB2X2

MACRO AOI2BB2X1
    CLASS CORE ;
    FOREIGN AOI2BB2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI2BB2XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.150 0.690 3.450 0.930 ;
        RECT  3.450 0.690 3.690 1.100 ;
        RECT  3.500 4.060 3.760 4.330 ;
        RECT  3.760 4.060 3.970 4.320 ;
        RECT  3.970 3.800 4.030 4.320 ;
        RECT  3.690 0.860 4.030 1.100 ;
        RECT  4.030 0.860 4.270 4.320 ;
        RECT  4.270 3.760 4.290 4.320 ;
        RECT  4.290 3.760 4.370 4.200 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.090 1.820 2.190 2.100 ;
        RECT  2.190 1.820 2.430 2.430 ;
        RECT  2.430 1.820 2.530 2.100 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.750 2.380 2.980 2.660 ;
        RECT  2.980 2.110 3.220 2.660 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.500 0.530 2.090 ;
        RECT  0.530 1.670 0.590 2.070 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.250 1.300 2.670 ;
        END
    END A0N
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 2.650 5.440 ;
        RECT  2.650 4.000 2.660 5.440 ;
        RECT  2.660 3.800 3.060 5.440 ;
        RECT  3.060 4.000 3.070 5.440 ;
        RECT  3.070 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 1.010 ;
        RECT  0.170 -0.400 0.570 1.130 ;
        RECT  0.570 -0.400 0.580 1.010 ;
        RECT  0.580 -0.400 1.930 0.400 ;
        RECT  1.930 -0.400 2.330 0.870 ;
        RECT  2.330 -0.400 3.970 0.400 ;
        RECT  3.970 -0.400 4.370 0.560 ;
        RECT  4.370 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.040 1.460 3.750 1.700 ;
        RECT  2.330 3.200 3.730 3.440 ;
        RECT  2.800 1.310 3.040 1.700 ;
        RECT  1.810 1.310 2.800 1.550 ;
        RECT  2.090 3.120 2.330 3.520 ;
        RECT  1.630 1.310 1.810 3.310 ;
        RECT  1.570 1.310 1.630 3.470 ;
        RECT  1.370 1.310 1.570 1.550 ;
        RECT  1.230 3.070 1.570 3.470 ;
        RECT  1.130 0.960 1.370 1.550 ;
    END
END AOI2BB2X1

MACRO AOI2BB1XL
    CLASS CORE ;
    FOREIGN AOI2BB1XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.130 1.150 2.770 1.390 ;
        RECT  2.770 1.150 3.010 4.000 ;
        RECT  3.010 3.510 3.090 4.000 ;
        RECT  3.090 3.510 3.100 3.770 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.430 2.760 1.930 3.220 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.820 1.330 2.250 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.620 0.550 3.220 ;
        RECT  0.550 2.810 0.620 3.210 ;
        END
    END A0N
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.420 5.440 ;
        RECT  1.420 4.480 1.820 5.440 ;
        RECT  1.820 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        RECT  0.940 -0.400 1.340 0.560 ;
        RECT  1.340 -0.400 2.740 0.400 ;
        RECT  2.740 -0.400 3.140 0.560 ;
        RECT  3.140 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.440 2.070 2.490 2.470 ;
        RECT  2.200 2.070 2.440 3.730 ;
        RECT  1.850 2.070 2.200 2.310 ;
        RECT  0.180 3.490 2.200 3.730 ;
        RECT  1.610 1.300 1.850 2.310 ;
        RECT  0.450 1.300 1.610 1.540 ;
    END
END AOI2BB1XL

MACRO AOI2BB1X4
    CLASS CORE ;
    FOREIGN AOI2BB1X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI2BB1XL ;
    SIZE 7.260 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.770 2.790 4.170 4.120 ;
        RECT  4.020 1.140 4.260 1.540 ;
        RECT  4.260 1.220 4.950 1.460 ;
        RECT  4.950 1.220 5.310 1.540 ;
        RECT  4.170 2.790 5.610 3.190 ;
        RECT  5.310 1.140 5.710 1.540 ;
        RECT  5.610 2.790 5.850 3.220 ;
        RECT  5.850 2.530 6.050 3.220 ;
        RECT  6.050 2.530 6.390 4.340 ;
        RECT  5.710 1.220 6.390 1.460 ;
        RECT  6.390 1.220 6.490 4.340 ;
        RECT  6.490 1.220 6.630 3.650 ;
        RECT  6.630 2.510 6.710 3.650 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 1.830 2.930 2.090 ;
        RECT  2.930 1.700 3.230 2.350 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.260 2.160 0.500 3.740 ;
        RECT  0.500 3.500 2.090 3.740 ;
        RECT  2.090 1.790 2.330 3.740 ;
        RECT  2.330 2.950 2.440 3.210 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 0.870 2.090 ;
        RECT  0.870 1.830 1.210 2.700 ;
        RECT  1.210 2.300 1.290 2.700 ;
        END
    END A0N
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 2.500 5.440 ;
        RECT  2.500 4.140 2.510 5.440 ;
        RECT  2.510 4.020 2.910 5.440 ;
        RECT  2.910 4.140 2.920 5.440 ;
        RECT  2.920 4.640 5.100 5.440 ;
        RECT  5.100 3.940 5.110 5.440 ;
        RECT  5.110 3.460 5.510 5.440 ;
        RECT  5.510 3.940 5.520 5.440 ;
        RECT  5.520 4.640 7.260 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.220 0.400 ;
        RECT  1.220 -0.400 1.230 0.790 ;
        RECT  1.230 -0.400 1.630 0.990 ;
        RECT  1.630 -0.400 1.640 0.790 ;
        RECT  1.640 -0.400 3.280 0.400 ;
        RECT  3.280 -0.400 3.290 0.670 ;
        RECT  3.290 -0.400 3.690 0.870 ;
        RECT  3.690 -0.400 3.700 0.670 ;
        RECT  3.700 -0.400 4.620 0.400 ;
        RECT  4.620 -0.400 4.630 0.670 ;
        RECT  4.630 -0.400 5.030 0.870 ;
        RECT  5.030 -0.400 5.040 0.670 ;
        RECT  5.040 -0.400 5.950 0.400 ;
        RECT  5.950 -0.400 5.960 0.670 ;
        RECT  5.960 -0.400 6.360 0.870 ;
        RECT  6.360 -0.400 6.370 0.670 ;
        RECT  6.370 -0.400 7.260 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.570 1.820 5.730 2.220 ;
        RECT  5.330 1.820 5.570 2.500 ;
        RECT  3.740 2.260 5.330 2.500 ;
        RECT  3.500 1.190 3.740 2.500 ;
        RECT  2.410 1.190 3.500 1.430 ;
        RECT  2.010 1.110 2.410 1.510 ;
        RECT  1.810 1.270 2.010 1.510 ;
        RECT  1.570 1.270 1.810 3.220 ;
        RECT  0.850 1.270 1.570 1.510 ;
        RECT  1.230 2.980 1.570 3.220 ;
        RECT  0.450 1.110 0.850 1.510 ;
    END
END AOI2BB1X4

MACRO AOI2BB1X2
    CLASS CORE ;
    FOREIGN AOI2BB1X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI2BB1XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.650 3.100 2.750 3.500 ;
        RECT  2.450 0.920 2.850 1.320 ;
        RECT  2.750 3.100 3.190 3.770 ;
        RECT  3.190 3.100 4.210 3.340 ;
        RECT  2.850 1.080 4.210 1.320 ;
        RECT  4.210 1.080 4.450 3.340 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.210 1.780 2.450 2.180 ;
        RECT  2.450 1.820 3.690 2.100 ;
        RECT  3.690 1.820 3.930 2.710 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 1.120 3.210 ;
        RECT  1.120 2.950 1.210 3.190 ;
        RECT  1.210 2.310 1.450 3.190 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.820 0.500 2.600 ;
        END
    END A0N
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.370 5.440 ;
        RECT  1.370 4.480 1.770 5.440 ;
        RECT  1.770 4.640 3.920 5.440 ;
        RECT  3.920 3.820 3.930 5.440 ;
        RECT  3.930 3.620 4.330 5.440 ;
        RECT  4.330 3.820 4.340 5.440 ;
        RECT  4.340 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 1.410 ;
        RECT  0.570 -0.400 1.680 0.400 ;
        RECT  1.680 -0.400 1.690 1.300 ;
        RECT  1.690 -0.400 2.090 1.420 ;
        RECT  2.090 -0.400 2.100 1.300 ;
        RECT  2.100 -0.400 3.270 0.400 ;
        RECT  3.270 -0.400 3.670 0.560 ;
        RECT  3.670 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.890 2.380 3.290 2.720 ;
        RECT  1.970 2.480 2.890 2.720 ;
        RECT  1.730 1.790 1.970 3.900 ;
        RECT  1.330 1.790 1.730 2.030 ;
        RECT  0.170 3.660 1.730 3.900 ;
        RECT  0.930 1.140 1.330 2.030 ;
    END
END AOI2BB1X2

MACRO AOI2BB1X1
    CLASS CORE ;
    FOREIGN AOI2BB1X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI2BB1XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.210 1.090 2.450 1.490 ;
        RECT  2.550 4.100 2.720 4.340 ;
        RECT  2.450 1.250 2.720 1.490 ;
        RECT  2.720 1.250 2.960 4.340 ;
        RECT  2.960 4.070 3.090 4.340 ;
        RECT  3.090 4.070 3.100 4.330 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.350 2.870 1.920 3.290 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.820 1.320 2.240 ;
        RECT  1.320 1.830 1.350 2.230 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.610 0.460 3.210 ;
        RECT  0.460 2.610 0.550 3.020 ;
        RECT  0.550 2.620 0.810 3.020 ;
        END
    END A0N
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.240 5.440 ;
        RECT  1.240 4.480 1.640 5.440 ;
        RECT  1.640 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.940 0.400 ;
        RECT  0.940 -0.400 1.340 0.560 ;
        RECT  1.340 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.190 1.870 2.430 3.820 ;
        RECT  1.880 1.870 2.190 2.110 ;
        RECT  0.170 3.580 2.190 3.820 ;
        RECT  1.640 1.310 1.880 2.110 ;
        RECT  0.450 1.310 1.640 1.550 ;
    END
END AOI2BB1X1

MACRO AOI22XL
    CLASS CORE ;
    FOREIGN AOI22XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.450 0.910 1.850 1.310 ;
        RECT  1.850 0.980 1.870 1.310 ;
        RECT  2.410 2.920 2.570 3.320 ;
        RECT  2.570 2.420 2.810 3.320 ;
        RECT  1.870 1.070 3.500 1.310 ;
        RECT  2.810 2.420 3.510 2.660 ;
        RECT  3.500 1.070 3.510 1.530 ;
        RECT  3.510 1.070 3.750 2.660 ;
        RECT  3.750 1.270 3.760 1.530 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.270 0.240 1.530 ;
        RECT  0.240 1.270 0.460 1.930 ;
        RECT  0.460 1.290 0.480 1.930 ;
        RECT  0.480 1.530 0.880 1.930 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 1.120 2.790 ;
        RECT  1.120 2.400 1.610 2.790 ;
        RECT  1.610 2.430 1.620 2.790 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.420 1.600 2.580 2.000 ;
        RECT  2.580 1.600 2.820 2.070 ;
        RECT  2.820 1.830 2.840 2.070 ;
        RECT  2.840 1.830 3.100 2.090 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.530 2.090 ;
        RECT  1.530 1.590 2.090 2.090 ;
        RECT  2.090 1.780 2.100 2.090 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.840 5.440 ;
        RECT  0.840 4.480 1.240 5.440 ;
        RECT  1.240 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 0.790 ;
        RECT  0.170 -0.400 0.570 0.990 ;
        RECT  0.570 -0.400 0.580 0.790 ;
        RECT  0.580 -0.400 2.730 0.400 ;
        RECT  2.730 -0.400 3.130 0.560 ;
        RECT  3.130 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.170 3.300 3.570 3.840 ;
        RECT  2.050 3.600 3.170 3.840 ;
        RECT  1.650 3.300 2.050 3.840 ;
        RECT  0.570 3.380 1.650 3.620 ;
        RECT  0.170 3.300 0.570 3.700 ;
    END
END AOI22XL

MACRO AOI22X4
    CLASS CORE ;
    FOREIGN AOI22X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI22XL ;
    SIZE 11.220 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.460 1.140 1.470 1.560 ;
        RECT  1.470 0.990 1.870 1.560 ;
        RECT  1.870 1.140 3.620 1.560 ;
        RECT  3.620 0.990 4.330 1.560 ;
        RECT  5.930 3.900 6.130 4.300 ;
        RECT  4.330 1.140 6.260 1.560 ;
        RECT  6.260 0.980 6.880 1.560 ;
        RECT  6.880 1.140 8.920 1.560 ;
        RECT  8.920 0.990 9.570 1.560 ;
        RECT  9.570 1.140 10.010 1.560 ;
        RECT  6.130 3.890 10.440 4.310 ;
        RECT  10.010 1.140 10.440 2.660 ;
        RECT  10.440 1.140 10.450 4.310 ;
        RECT  10.450 1.960 10.860 4.310 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.420 1.820 3.380 2.230 ;
        RECT  3.380 1.820 4.860 2.100 ;
        RECT  4.860 1.820 5.260 2.220 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.020 2.270 1.420 2.670 ;
        RECT  1.420 2.380 1.670 2.750 ;
        RECT  1.670 2.390 1.780 2.750 ;
        RECT  1.780 2.510 3.800 2.750 ;
        RECT  3.800 2.390 4.200 2.790 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.630 2.500 5.790 2.740 ;
        RECT  5.790 1.840 6.200 2.740 ;
        RECT  6.200 1.840 7.460 2.080 ;
        RECT  7.460 1.830 7.720 2.090 ;
        RECT  7.720 1.840 8.350 2.080 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.440 2.400 6.710 2.640 ;
        RECT  6.710 2.380 9.280 2.660 ;
        RECT  9.280 2.260 9.680 2.660 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.240 5.440 ;
        RECT  1.240 4.060 1.250 5.440 ;
        RECT  1.250 3.580 1.650 5.440 ;
        RECT  1.650 4.060 1.660 5.440 ;
        RECT  1.660 4.640 2.800 5.440 ;
        RECT  2.800 4.060 2.810 5.440 ;
        RECT  2.810 3.580 3.210 5.440 ;
        RECT  3.210 4.060 3.220 5.440 ;
        RECT  3.220 4.640 4.360 5.440 ;
        RECT  4.360 4.060 4.370 5.440 ;
        RECT  4.370 3.580 4.770 5.440 ;
        RECT  4.770 4.060 4.780 5.440 ;
        RECT  4.780 4.640 11.220 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 2.690 0.400 ;
        RECT  2.690 -0.400 2.700 0.670 ;
        RECT  2.700 -0.400 3.100 0.870 ;
        RECT  3.100 -0.400 3.110 0.670 ;
        RECT  3.110 -0.400 5.140 0.400 ;
        RECT  5.140 -0.400 5.150 0.670 ;
        RECT  5.150 -0.400 5.550 0.870 ;
        RECT  5.550 -0.400 5.560 0.670 ;
        RECT  5.560 -0.400 7.580 0.400 ;
        RECT  7.580 -0.400 7.590 0.670 ;
        RECT  7.590 -0.400 7.990 0.870 ;
        RECT  7.990 -0.400 8.000 0.670 ;
        RECT  8.000 -0.400 11.220 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  9.770 3.070 10.170 3.610 ;
        RECT  8.670 3.070 9.770 3.310 ;
        RECT  8.270 3.070 8.670 3.620 ;
        RECT  7.110 3.070 8.270 3.310 ;
        RECT  6.710 3.070 7.110 3.610 ;
        RECT  5.550 3.070 6.710 3.310 ;
        RECT  5.150 3.070 5.550 3.610 ;
        RECT  3.990 3.070 5.150 3.310 ;
        RECT  3.590 3.070 3.990 3.610 ;
        RECT  2.430 3.070 3.590 3.310 ;
        RECT  2.030 3.070 2.430 3.610 ;
        RECT  0.930 3.070 2.030 3.310 ;
        RECT  0.530 3.070 0.930 3.610 ;
    END
END AOI22X4

MACRO AOI22X2
    CLASS CORE ;
    FOREIGN AOI22X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI22XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.050 0.670 2.260 0.910 ;
        RECT  2.260 0.670 2.500 1.180 ;
        RECT  4.090 3.180 5.480 3.420 ;
        RECT  5.480 2.940 5.800 3.420 ;
        RECT  2.500 0.940 6.050 1.180 ;
        RECT  5.800 2.940 6.190 3.200 ;
        RECT  6.050 0.940 6.190 1.390 ;
        RECT  6.190 0.940 6.430 3.200 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.070 1.500 1.270 1.900 ;
        RECT  1.270 1.490 1.430 1.910 ;
        RECT  1.430 1.270 1.870 1.910 ;
        RECT  1.870 1.490 3.230 1.910 ;
        RECT  3.230 1.500 3.430 1.900 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.680 2.330 2.330 2.730 ;
        RECT  2.330 2.320 2.590 2.740 ;
        RECT  2.590 2.330 2.640 2.730 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 2.390 3.650 2.650 ;
        RECT  3.650 2.350 4.050 2.750 ;
        RECT  4.050 2.350 4.320 2.670 ;
        RECT  4.320 2.430 5.670 2.670 ;
        RECT  5.670 2.240 5.910 2.670 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.340 1.830 5.170 2.100 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.280 5.440 ;
        RECT  1.280 3.980 1.290 5.440 ;
        RECT  1.290 3.780 1.690 5.440 ;
        RECT  1.690 3.980 1.700 5.440 ;
        RECT  1.700 4.640 2.620 5.440 ;
        RECT  2.620 3.980 2.630 5.440 ;
        RECT  2.630 3.780 3.030 5.440 ;
        RECT  3.030 3.980 3.040 5.440 ;
        RECT  3.040 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.820 0.400 ;
        RECT  0.820 -0.400 0.830 0.790 ;
        RECT  0.830 -0.400 1.230 0.990 ;
        RECT  1.230 -0.400 1.240 0.790 ;
        RECT  1.240 -0.400 3.330 0.400 ;
        RECT  3.330 -0.400 3.730 0.560 ;
        RECT  3.730 -0.400 5.490 0.400 ;
        RECT  5.490 -0.400 6.300 0.560 ;
        RECT  6.300 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.700 3.780 6.420 4.180 ;
        RECT  3.300 3.100 3.700 4.180 ;
        RECT  2.360 3.180 3.300 3.420 ;
        RECT  1.960 3.100 2.360 3.500 ;
        RECT  1.070 3.180 1.960 3.420 ;
        RECT  0.670 3.100 1.070 3.500 ;
    END
END AOI22X2

MACRO AOI22X1
    CLASS CORE ;
    FOREIGN AOI22X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI22XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.390 0.670 2.150 0.910 ;
        RECT  2.150 0.670 2.390 1.340 ;
        RECT  2.390 0.960 2.430 1.340 ;
        RECT  2.560 2.830 2.960 3.230 ;
        RECT  2.960 2.830 3.410 3.070 ;
        RECT  2.430 1.100 3.500 1.340 ;
        RECT  3.410 2.660 3.510 3.070 ;
        RECT  3.500 1.100 3.510 1.530 ;
        RECT  3.510 1.100 3.740 3.070 ;
        RECT  3.740 1.270 3.750 3.070 ;
        RECT  3.750 1.270 3.760 1.530 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.270 0.460 1.890 ;
        RECT  0.460 1.490 0.740 1.890 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.250 1.220 2.670 ;
        RECT  1.220 2.260 1.610 2.660 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.760 1.580 3.140 2.220 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.270 1.630 1.530 ;
        RECT  1.630 1.270 1.780 1.860 ;
        RECT  1.780 1.290 1.870 1.860 ;
        RECT  1.870 1.620 2.060 1.860 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.920 5.440 ;
        RECT  0.920 4.480 1.320 5.440 ;
        RECT  1.320 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 0.780 ;
        RECT  0.170 -0.400 0.570 0.900 ;
        RECT  0.570 -0.400 0.580 0.780 ;
        RECT  0.580 -0.400 2.670 0.400 ;
        RECT  2.670 -0.400 3.070 0.560 ;
        RECT  3.070 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.520 3.570 3.720 3.970 ;
        RECT  0.370 3.560 3.520 3.980 ;
        RECT  0.170 3.570 0.370 3.970 ;
    END
END AOI22X1

MACRO AOI222XL
    CLASS CORE ;
    FOREIGN AOI222XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.170 0.670 0.850 0.910 ;
        RECT  0.850 0.670 1.090 1.340 ;
        RECT  1.090 0.960 1.110 1.340 ;
        RECT  1.110 1.100 2.670 1.340 ;
        RECT  2.670 0.980 2.830 1.340 ;
        RECT  2.830 0.750 2.910 1.340 ;
        RECT  2.910 0.750 3.070 1.220 ;
        RECT  3.070 0.750 4.120 0.990 ;
        RECT  4.120 0.750 4.360 1.550 ;
        RECT  4.010 2.850 4.730 3.090 ;
        RECT  4.730 2.410 4.820 3.090 ;
        RECT  4.820 2.390 4.830 3.090 ;
        RECT  4.360 1.310 4.830 1.550 ;
        RECT  4.830 1.310 4.970 3.090 ;
        RECT  4.970 1.310 5.070 2.650 ;
        RECT  5.070 2.390 5.080 2.650 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.630 1.300 2.100 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.160 1.210 0.500 1.860 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.390 1.700 2.650 ;
        RECT  1.700 1.720 1.780 2.650 ;
        RECT  1.780 1.720 2.100 2.640 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.420 1.630 2.580 2.030 ;
        RECT  2.580 1.630 2.820 2.070 ;
        RECT  2.820 1.830 2.840 2.070 ;
        RECT  2.840 1.830 3.100 2.090 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 1.830 4.220 2.090 ;
        RECT  4.220 1.830 4.420 2.570 ;
        RECT  4.420 1.840 4.460 2.570 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.450 1.260 3.760 1.880 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 0.250 5.440 ;
        RECT  0.250 4.460 1.090 5.440 ;
        RECT  1.090 4.480 1.170 5.440 ;
        RECT  1.170 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.380 0.400 ;
        RECT  1.380 -0.400 1.390 0.690 ;
        RECT  1.390 -0.400 1.790 0.810 ;
        RECT  1.790 -0.400 1.800 0.690 ;
        RECT  1.800 -0.400 4.640 0.400 ;
        RECT  4.640 -0.400 5.040 0.560 ;
        RECT  5.040 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.150 4.130 5.000 4.370 ;
        RECT  2.630 2.770 3.030 3.170 ;
        RECT  1.150 2.930 2.630 3.170 ;
        RECT  0.750 2.800 1.150 3.200 ;
    END
END AOI222XL

MACRO AOI222X4
    CLASS CORE ;
    FOREIGN AOI222X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI222XL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.710 2.380 7.000 3.780 ;
        RECT  6.600 1.300 7.000 1.540 ;
        RECT  7.000 1.300 7.150 3.780 ;
        RECT  7.150 2.990 7.230 3.650 ;
        RECT  7.150 1.300 7.240 2.620 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.150 1.530 0.510 2.090 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.680 1.210 2.100 ;
        RECT  1.210 1.690 1.550 2.100 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.380 2.080 2.660 ;
        RECT  2.080 2.250 2.440 2.660 ;
        RECT  2.440 2.250 2.480 2.650 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.800 1.670 3.260 2.090 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 1.080 4.640 1.540 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.410 2.380 3.680 2.660 ;
        RECT  3.680 2.340 3.850 2.660 ;
        RECT  3.850 2.340 4.080 2.640 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 5.930 5.440 ;
        RECT  5.930 4.630 6.030 5.440 ;
        RECT  6.030 3.770 6.450 5.440 ;
        RECT  6.450 4.640 7.540 5.440 ;
        RECT  7.540 4.250 7.550 5.440 ;
        RECT  7.550 4.050 7.950 5.440 ;
        RECT  7.950 4.250 7.960 5.440 ;
        RECT  7.960 4.640 8.580 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 1.260 ;
        RECT  0.570 -0.400 0.700 0.410 ;
        RECT  0.700 -0.400 2.130 0.400 ;
        RECT  2.130 -0.400 2.530 0.560 ;
        RECT  2.530 -0.400 4.470 0.400 ;
        RECT  4.470 -0.400 4.870 0.790 ;
        RECT  4.870 -0.400 5.980 0.400 ;
        RECT  5.980 -0.400 5.990 0.740 ;
        RECT  5.990 -0.400 6.390 0.940 ;
        RECT  6.390 -0.400 6.400 0.740 ;
        RECT  6.400 -0.400 7.240 0.400 ;
        RECT  7.240 -0.400 7.250 0.740 ;
        RECT  7.250 -0.400 7.650 0.940 ;
        RECT  7.650 -0.400 7.660 0.740 ;
        RECT  7.660 -0.400 8.580 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.320 1.870 6.760 2.110 ;
        RECT  6.080 1.410 6.320 3.100 ;
        RECT  5.590 1.410 6.080 1.650 ;
        RECT  5.830 2.860 6.080 3.100 ;
        RECT  5.430 2.860 5.830 3.260 ;
        RECT  4.600 2.340 5.800 2.580 ;
        RECT  5.190 1.250 5.590 1.650 ;
        RECT  2.080 4.130 5.100 4.370 ;
        RECT  4.360 1.810 4.600 3.340 ;
        RECT  3.790 1.810 4.360 2.050 ;
        RECT  4.110 2.940 4.360 3.340 ;
        RECT  3.550 1.060 3.790 2.050 ;
        RECT  3.190 1.060 3.550 1.380 ;
        RECT  1.790 1.060 3.190 1.300 ;
        RECT  2.670 3.040 3.070 3.440 ;
        RECT  1.070 3.040 2.670 3.280 ;
        RECT  1.390 0.900 1.790 1.300 ;
        RECT  0.830 3.040 1.070 3.440 ;
    END
END AOI222X4

MACRO AOI222X2
    CLASS CORE ;
    FOREIGN AOI222X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI222XL ;
    SIZE 9.900 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.390 1.030 1.790 1.430 ;
        RECT  1.790 1.190 4.630 1.430 ;
        RECT  4.630 0.810 5.030 1.430 ;
        RECT  5.030 0.960 5.170 1.430 ;
        RECT  5.170 1.190 7.070 1.430 ;
        RECT  6.790 2.940 7.190 3.340 ;
        RECT  7.070 0.810 7.470 1.430 ;
        RECT  7.190 2.940 7.610 3.260 ;
        RECT  7.610 3.020 8.120 3.260 ;
        RECT  8.120 2.950 8.130 3.260 ;
        RECT  8.130 2.940 8.280 3.340 ;
        RECT  7.470 1.190 8.370 1.430 ;
        RECT  8.370 1.190 8.470 1.520 ;
        RECT  8.280 2.790 8.530 3.340 ;
        RECT  8.530 2.790 8.660 3.260 ;
        RECT  8.470 1.190 8.660 1.540 ;
        RECT  8.660 1.190 8.900 3.260 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.460 2.250 0.860 2.650 ;
        RECT  0.860 2.390 1.120 2.650 ;
        RECT  1.120 2.400 2.770 2.640 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.350 1.760 1.930 2.100 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.670 2.090 ;
        RECT  3.670 1.710 4.310 2.110 ;
        RECT  4.310 1.850 5.170 2.090 ;
        RECT  5.170 1.850 5.380 2.100 ;
        RECT  5.380 1.850 5.780 2.320 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 2.390 4.420 2.650 ;
        RECT  4.420 2.400 5.060 2.640 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.110 1.840 6.140 2.080 ;
        RECT  6.140 1.830 6.400 2.090 ;
        RECT  6.400 1.840 8.130 2.080 ;
        RECT  8.130 1.840 8.370 2.320 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.800 2.390 7.050 2.650 ;
        RECT  7.050 2.380 7.740 2.660 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.000 0.170 5.440 ;
        RECT  0.170 3.800 0.570 5.440 ;
        RECT  0.570 4.000 0.580 5.440 ;
        RECT  0.580 4.640 1.450 5.440 ;
        RECT  1.450 4.000 1.460 5.440 ;
        RECT  1.460 3.800 1.860 5.440 ;
        RECT  1.860 4.000 1.870 5.440 ;
        RECT  1.870 4.640 2.740 5.440 ;
        RECT  2.740 4.000 2.750 5.440 ;
        RECT  2.750 3.800 3.150 5.440 ;
        RECT  3.150 4.000 3.160 5.440 ;
        RECT  3.160 4.640 9.900 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.180 0.400 ;
        RECT  0.180 -0.400 0.190 1.230 ;
        RECT  0.190 -0.400 0.590 1.430 ;
        RECT  0.590 -0.400 0.600 1.230 ;
        RECT  0.600 -0.400 2.660 0.400 ;
        RECT  2.660 -0.400 2.670 0.710 ;
        RECT  2.670 -0.400 3.070 0.910 ;
        RECT  3.070 -0.400 3.080 0.710 ;
        RECT  3.080 -0.400 3.400 0.400 ;
        RECT  3.400 -0.400 3.410 0.710 ;
        RECT  3.410 -0.400 3.810 0.910 ;
        RECT  3.810 -0.400 3.820 0.710 ;
        RECT  3.820 -0.400 5.840 0.400 ;
        RECT  5.840 -0.400 5.850 0.700 ;
        RECT  5.850 -0.400 6.250 0.900 ;
        RECT  6.250 -0.400 6.260 0.700 ;
        RECT  6.260 -0.400 8.260 0.400 ;
        RECT  8.260 -0.400 8.270 0.700 ;
        RECT  8.270 -0.400 8.670 0.900 ;
        RECT  8.670 -0.400 8.680 0.700 ;
        RECT  8.680 -0.400 9.900 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  8.950 3.800 9.150 4.200 ;
        RECT  3.690 3.790 8.950 4.210 ;
        RECT  5.450 2.940 5.850 3.340 ;
        RECT  4.510 3.020 5.450 3.260 ;
        RECT  4.110 2.940 4.510 3.340 ;
        RECT  2.530 3.020 4.110 3.260 ;
        RECT  3.490 3.800 3.690 4.200 ;
        RECT  2.130 2.940 2.530 3.340 ;
        RECT  1.190 3.020 2.130 3.260 ;
        RECT  0.790 2.940 1.190 3.340 ;
    END
END AOI222X2

MACRO AOI222X1
    CLASS CORE ;
    FOREIGN AOI222X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI222XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.170 1.030 0.570 1.430 ;
        RECT  0.570 1.030 2.090 1.270 ;
        RECT  2.090 0.980 2.140 1.270 ;
        RECT  2.140 0.750 2.380 1.270 ;
        RECT  2.380 0.750 3.460 0.990 ;
        RECT  3.460 0.750 3.700 1.100 ;
        RECT  4.110 2.930 4.510 3.330 ;
        RECT  4.510 2.930 4.730 3.220 ;
        RECT  4.730 2.930 4.830 3.200 ;
        RECT  3.700 0.860 5.390 1.100 ;
        RECT  4.830 2.930 5.490 3.170 ;
        RECT  5.480 2.390 5.490 2.650 ;
        RECT  5.390 0.860 5.490 1.260 ;
        RECT  5.490 0.860 5.730 3.170 ;
        RECT  5.730 2.390 5.740 2.650 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.100 2.340 1.650 2.660 ;
        RECT  1.650 2.380 1.870 2.660 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.290 2.090 ;
        RECT  0.290 1.830 0.460 2.580 ;
        RECT  0.460 1.850 0.530 2.580 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.110 1.850 2.180 2.550 ;
        RECT  2.180 1.830 2.350 2.550 ;
        RECT  2.350 1.830 2.440 2.090 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.770 1.270 3.140 1.800 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.360 1.450 5.080 2.090 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.510 1.900 3.750 2.620 ;
        RECT  3.750 2.380 4.160 2.620 ;
        RECT  4.160 2.380 4.410 2.650 ;
        RECT  4.410 2.390 4.420 2.650 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.990 0.170 5.440 ;
        RECT  0.170 3.790 0.570 5.440 ;
        RECT  0.570 3.990 0.580 5.440 ;
        RECT  0.580 4.640 1.400 5.440 ;
        RECT  1.400 3.990 1.410 5.440 ;
        RECT  1.410 3.790 1.810 5.440 ;
        RECT  1.810 3.990 1.820 5.440 ;
        RECT  1.820 4.630 2.000 5.440 ;
        RECT  2.000 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.450 0.400 ;
        RECT  1.450 -0.400 1.850 0.560 ;
        RECT  1.850 -0.400 4.200 0.400 ;
        RECT  4.200 -0.400 4.600 0.560 ;
        RECT  4.600 -0.400 5.940 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.930 3.790 5.130 4.190 ;
        RECT  2.350 3.780 4.930 4.200 ;
        RECT  2.770 2.930 3.170 3.330 ;
        RECT  1.110 2.990 2.770 3.230 ;
        RECT  2.150 3.790 2.350 4.190 ;
        RECT  0.870 2.910 1.110 3.310 ;
    END
END AOI222X1

MACRO AOI221XL
    CLASS CORE ;
    FOREIGN AOI221XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.390 0.670 1.770 0.910 ;
        RECT  1.770 0.670 1.900 0.980 ;
        RECT  1.900 0.670 2.140 1.100 ;
        RECT  2.140 0.720 2.190 1.100 ;
        RECT  2.190 0.860 3.590 1.100 ;
        RECT  3.590 0.860 3.600 1.260 ;
        RECT  3.600 0.840 4.000 1.260 ;
        RECT  4.120 2.500 4.160 3.170 ;
        RECT  4.160 2.390 4.170 3.170 ;
        RECT  4.000 1.010 4.170 1.260 ;
        RECT  4.170 1.010 4.410 3.170 ;
        RECT  4.410 2.390 4.420 2.650 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.460 1.650 3.500 2.640 ;
        RECT  3.500 1.650 3.700 2.650 ;
        RECT  3.700 2.390 3.760 2.650 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.490 0.500 2.090 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 1.340 2.890 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.480 1.540 2.720 2.070 ;
        RECT  2.720 1.820 2.750 2.070 ;
        RECT  2.750 1.830 2.840 2.070 ;
        RECT  2.840 1.830 3.100 2.090 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.730 2.090 ;
        RECT  1.730 1.830 1.780 2.380 ;
        RECT  1.780 1.840 1.970 2.380 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.320 5.440 ;
        RECT  1.320 4.480 1.720 5.440 ;
        RECT  1.720 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.250 0.400 ;
        RECT  0.250 -0.400 0.490 0.890 ;
        RECT  0.490 -0.400 2.710 0.400 ;
        RECT  2.710 -0.400 3.110 0.560 ;
        RECT  3.110 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.050 4.130 3.580 4.370 ;
        RECT  2.680 2.770 2.920 3.420 ;
        RECT  0.740 3.180 2.680 3.420 ;
    END
END AOI221XL

MACRO AOI221X4
    CLASS CORE ;
    FOREIGN AOI221X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI221XL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  6.590 1.000 6.710 1.400 ;
        RECT  6.590 3.210 6.720 4.190 ;
        RECT  6.710 1.000 6.720 2.660 ;
        RECT  6.720 1.000 6.990 4.190 ;
        RECT  6.990 1.000 7.000 3.240 ;
        RECT  7.000 1.000 7.050 2.660 ;
        RECT  7.050 1.260 7.150 2.660 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.820 3.760 2.090 ;
        RECT  3.760 1.820 4.060 2.080 ;
        RECT  4.060 1.630 4.300 2.080 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.460 2.650 ;
        RECT  0.460 2.390 0.530 2.630 ;
        RECT  0.530 1.970 0.770 2.630 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 1.010 3.210 ;
        RECT  1.010 2.490 1.120 3.210 ;
        RECT  1.120 2.490 1.250 3.200 ;
        RECT  1.250 2.490 1.530 2.730 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.780 2.060 3.140 2.650 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.780 2.090 ;
        RECT  1.780 1.830 1.840 2.080 ;
        RECT  1.840 1.680 2.240 2.080 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 4.480 0.560 5.440 ;
        RECT  0.560 4.640 1.490 5.440 ;
        RECT  1.490 4.480 1.890 5.440 ;
        RECT  1.890 4.640 5.820 5.440 ;
        RECT  5.820 3.730 5.830 5.440 ;
        RECT  5.830 3.240 6.230 5.440 ;
        RECT  6.230 3.730 6.240 5.440 ;
        RECT  6.240 4.640 7.340 5.440 ;
        RECT  7.340 3.700 7.350 5.440 ;
        RECT  7.350 3.210 7.750 5.440 ;
        RECT  7.750 3.700 7.760 5.440 ;
        RECT  7.760 4.640 7.920 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.380 0.400 ;
        RECT  0.380 -0.400 0.780 1.450 ;
        RECT  0.780 -0.400 2.880 0.400 ;
        RECT  2.880 -0.400 3.280 0.560 ;
        RECT  3.280 -0.400 5.820 0.400 ;
        RECT  5.820 -0.400 5.830 1.030 ;
        RECT  5.830 -0.400 6.230 1.230 ;
        RECT  6.230 -0.400 6.240 1.030 ;
        RECT  6.240 -0.400 7.340 0.400 ;
        RECT  7.340 -0.400 7.350 0.670 ;
        RECT  7.350 -0.400 7.750 0.870 ;
        RECT  7.750 -0.400 7.760 0.670 ;
        RECT  7.760 -0.400 7.920 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.230 2.050 6.470 2.450 ;
        RECT  5.550 2.210 6.230 2.450 ;
        RECT  5.470 1.120 5.550 4.200 ;
        RECT  5.310 1.120 5.470 4.210 ;
        RECT  5.150 1.120 5.310 1.520 ;
        RECT  5.070 3.810 5.310 4.210 ;
        RECT  4.870 2.050 5.030 2.450 ;
        RECT  4.870 3.060 4.950 3.460 ;
        RECT  4.630 1.050 4.870 3.460 ;
        RECT  2.590 1.050 4.630 1.290 ;
        RECT  4.550 3.060 4.630 3.460 ;
        RECT  3.740 3.480 4.140 3.900 ;
        RECT  2.620 3.660 3.740 3.900 ;
        RECT  2.980 3.030 3.380 3.380 ;
        RECT  1.890 3.030 2.980 3.270 ;
        RECT  2.220 3.560 2.620 3.900 ;
        RECT  2.350 1.050 2.590 1.370 ;
        RECT  1.600 1.130 2.350 1.370 ;
        RECT  1.650 3.030 1.890 3.730 ;
        RECT  0.880 3.490 1.650 3.730 ;
    END
END AOI221X4

MACRO AOI221X2
    CLASS CORE ;
    FOREIGN AOI221X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI221XL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.490 0.760 2.360 1.000 ;
        RECT  2.360 0.760 2.600 1.530 ;
        RECT  2.600 1.260 2.750 1.530 ;
        RECT  2.750 1.280 2.850 1.530 ;
        RECT  2.850 1.290 3.560 1.530 ;
        RECT  3.560 0.750 3.800 1.530 ;
        RECT  3.800 0.750 5.010 0.990 ;
        RECT  5.010 0.750 5.250 1.180 ;
        RECT  5.250 0.940 6.540 1.180 ;
        RECT  6.800 2.950 6.810 3.210 ;
        RECT  6.810 2.870 6.850 3.210 ;
        RECT  6.540 0.940 6.940 1.350 ;
        RECT  6.940 1.110 7.050 1.350 ;
        RECT  6.850 2.870 7.250 3.290 ;
        RECT  7.050 1.110 7.250 1.540 ;
        RECT  7.250 1.110 7.490 3.110 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.480 1.830 5.740 2.090 ;
        RECT  5.740 1.840 6.490 2.080 ;
        RECT  6.490 1.820 6.570 2.100 ;
        RECT  6.570 1.800 6.970 2.200 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.510 2.200 2.180 2.440 ;
        RECT  2.180 2.200 2.440 2.650 ;
        RECT  2.440 2.200 2.770 2.440 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.270 1.120 1.530 ;
        RECT  1.120 1.280 1.520 1.520 ;
        RECT  1.520 1.280 1.920 1.790 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 1.830 3.650 2.090 ;
        RECT  3.650 1.830 3.760 2.610 ;
        RECT  3.760 1.840 3.890 2.610 ;
        RECT  3.890 2.370 6.050 2.610 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.160 1.270 4.170 1.530 ;
        RECT  4.170 1.270 4.500 1.700 ;
        RECT  4.500 1.460 5.130 1.700 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.940 0.170 5.440 ;
        RECT  0.170 3.740 0.570 5.440 ;
        RECT  0.570 3.940 0.580 5.440 ;
        RECT  0.580 4.640 1.460 5.440 ;
        RECT  1.460 3.940 1.470 5.440 ;
        RECT  1.470 3.740 1.870 5.440 ;
        RECT  1.870 3.940 1.880 5.440 ;
        RECT  1.880 4.640 2.760 5.440 ;
        RECT  2.760 3.940 2.770 5.440 ;
        RECT  2.770 3.740 3.170 5.440 ;
        RECT  3.170 3.940 3.180 5.440 ;
        RECT  3.180 4.640 8.580 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.260 0.400 ;
        RECT  0.260 -0.400 0.270 0.790 ;
        RECT  0.270 -0.400 0.670 0.990 ;
        RECT  0.670 -0.400 0.680 0.790 ;
        RECT  0.680 -0.400 2.870 0.400 ;
        RECT  2.870 -0.400 2.880 0.810 ;
        RECT  2.880 -0.400 3.280 1.010 ;
        RECT  3.280 -0.400 3.290 0.810 ;
        RECT  3.290 -0.400 5.740 0.400 ;
        RECT  5.740 -0.400 6.140 0.560 ;
        RECT  6.140 -0.400 8.580 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  7.670 3.740 7.870 4.140 ;
        RECT  3.710 3.730 7.670 4.150 ;
        RECT  5.490 2.890 5.890 3.290 ;
        RECT  4.530 2.970 5.490 3.210 ;
        RECT  4.130 2.890 4.530 3.290 ;
        RECT  1.190 2.950 4.130 3.190 ;
        RECT  3.510 3.740 3.710 4.140 ;
        RECT  0.790 2.890 1.190 3.290 ;
    END
END AOI221X2

MACRO AOI221X1
    CLASS CORE ;
    FOREIGN AOI221X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI221XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.390 0.670 2.200 0.910 ;
        RECT  2.200 0.670 2.440 1.190 ;
        RECT  2.440 0.950 3.620 1.190 ;
        RECT  4.140 2.640 4.170 3.230 ;
        RECT  3.620 0.870 4.170 1.270 ;
        RECT  4.170 0.870 4.300 3.230 ;
        RECT  4.300 1.030 4.410 3.230 ;
        RECT  4.410 2.640 4.450 3.230 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 2.390 3.560 2.650 ;
        RECT  3.560 1.550 3.760 2.650 ;
        RECT  3.760 1.550 3.800 2.640 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.180 1.270 0.510 1.860 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 0.970 2.090 ;
        RECT  0.970 1.830 1.120 2.420 ;
        RECT  1.120 1.850 1.210 2.420 ;
        RECT  1.210 2.180 1.430 2.420 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.370 1.640 2.840 1.880 ;
        RECT  2.840 1.640 3.090 2.090 ;
        RECT  3.090 1.830 3.100 2.090 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.260 1.930 1.790 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.890 0.170 5.440 ;
        RECT  0.170 3.690 0.570 5.440 ;
        RECT  0.570 3.890 0.580 5.440 ;
        RECT  0.580 4.640 1.400 5.440 ;
        RECT  1.400 3.890 1.410 5.440 ;
        RECT  1.410 3.690 1.810 5.440 ;
        RECT  1.810 3.890 1.820 5.440 ;
        RECT  1.820 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 0.670 ;
        RECT  0.170 -0.400 0.570 0.790 ;
        RECT  0.570 -0.400 0.580 0.670 ;
        RECT  0.580 -0.400 2.760 0.400 ;
        RECT  2.760 -0.400 3.160 0.560 ;
        RECT  3.160 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.840 3.550 3.850 3.970 ;
        RECT  3.440 3.550 3.840 4.090 ;
        RECT  2.350 3.550 3.440 3.970 ;
        RECT  1.110 2.900 3.170 3.140 ;
        RECT  2.150 3.560 2.350 3.960 ;
        RECT  0.870 2.820 1.110 3.220 ;
    END
END AOI221X1

MACRO AOI21XL
    CLASS CORE ;
    FOREIGN AOI21XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.390 1.090 1.790 1.490 ;
        RECT  2.450 3.220 2.550 3.620 ;
        RECT  2.550 3.220 2.850 3.630 ;
        RECT  2.840 2.390 2.850 2.650 ;
        RECT  1.790 1.250 2.850 1.490 ;
        RECT  2.850 1.250 3.090 3.630 ;
        RECT  3.090 2.390 3.100 3.630 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.950 1.610 3.210 ;
        RECT  1.610 2.940 1.870 3.210 ;
        RECT  1.870 2.940 1.880 3.200 ;
        RECT  1.880 2.350 2.140 3.200 ;
        RECT  2.140 2.350 2.280 2.750 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.950 0.210 3.210 ;
        RECT  0.210 1.900 0.330 3.210 ;
        RECT  0.330 1.740 0.450 3.210 ;
        RECT  0.450 2.950 0.460 3.210 ;
        RECT  0.450 1.740 0.730 2.140 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 0.970 2.650 ;
        RECT  0.970 1.840 1.120 2.650 ;
        RECT  1.120 1.840 1.210 2.630 ;
        RECT  1.210 1.840 1.550 2.080 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.780 5.440 ;
        RECT  0.780 4.480 1.180 5.440 ;
        RECT  1.180 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 1.490 ;
        RECT  0.570 -0.400 2.160 0.400 ;
        RECT  2.160 -0.400 2.560 0.560 ;
        RECT  2.560 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  0.170 3.490 2.050 3.730 ;
    END
END AOI21XL

MACRO AOI21X4
    CLASS CORE ;
    FOREIGN AOI21X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI21XL ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.830 1.070 1.030 1.470 ;
        RECT  1.030 1.060 1.430 1.480 ;
        RECT  1.430 0.700 1.870 2.100 ;
        RECT  1.870 1.150 3.280 1.470 ;
        RECT  3.280 1.060 3.680 1.470 ;
        RECT  3.680 1.150 4.950 1.470 ;
        RECT  4.950 1.150 5.270 1.540 ;
        RECT  5.270 1.140 5.470 1.540 ;
        RECT  5.600 3.630 5.610 4.050 ;
        RECT  5.610 3.480 6.010 4.050 ;
        RECT  6.010 3.630 7.010 4.050 ;
        RECT  7.010 3.630 7.050 4.200 ;
        RECT  5.470 1.130 7.050 1.550 ;
        RECT  7.050 1.130 7.470 4.210 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.290 1.820 6.790 2.220 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.140 1.740 2.540 2.080 ;
        RECT  2.540 1.740 4.160 1.980 ;
        RECT  4.160 1.740 4.350 2.090 ;
        RECT  4.350 1.740 4.590 2.380 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.920 1.750 1.160 2.650 ;
        RECT  1.160 2.410 2.960 2.650 ;
        RECT  2.960 2.260 3.750 2.650 ;
        RECT  3.750 2.390 3.760 2.650 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.920 5.440 ;
        RECT  0.920 3.680 0.930 5.440 ;
        RECT  0.930 3.480 1.330 5.440 ;
        RECT  1.330 3.680 1.340 5.440 ;
        RECT  1.340 4.640 2.480 5.440 ;
        RECT  2.480 3.680 2.490 5.440 ;
        RECT  2.490 3.480 2.890 5.440 ;
        RECT  2.890 3.680 2.900 5.440 ;
        RECT  2.900 4.640 4.040 5.440 ;
        RECT  4.040 3.680 4.050 5.440 ;
        RECT  4.050 3.480 4.450 5.440 ;
        RECT  4.450 3.680 4.460 5.440 ;
        RECT  4.460 4.640 7.920 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 2.140 0.400 ;
        RECT  2.140 -0.400 2.380 0.870 ;
        RECT  2.380 -0.400 4.570 0.400 ;
        RECT  4.570 -0.400 4.970 0.560 ;
        RECT  4.970 -0.400 5.970 0.400 ;
        RECT  5.970 -0.400 6.370 0.560 ;
        RECT  6.370 -0.400 7.920 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.380 2.960 6.780 3.360 ;
        RECT  5.220 2.960 6.380 3.200 ;
        RECT  4.820 2.960 5.220 3.360 ;
        RECT  3.670 2.960 4.820 3.200 ;
        RECT  3.270 2.960 3.670 3.360 ;
        RECT  2.100 2.960 3.270 3.200 ;
        RECT  1.700 2.960 2.100 3.360 ;
        RECT  0.610 2.960 1.700 3.200 ;
        RECT  0.210 2.960 0.610 3.360 ;
    END
END AOI21X4

MACRO AOI21X2
    CLASS CORE ;
    FOREIGN AOI21X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI21XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.190 0.750 0.830 0.990 ;
        RECT  0.830 0.750 1.070 1.430 ;
        RECT  1.070 0.960 1.110 1.430 ;
        RECT  1.110 1.190 2.430 1.430 ;
        RECT  2.430 1.190 2.910 1.520 ;
        RECT  3.610 2.970 3.770 3.370 ;
        RECT  2.910 1.280 3.770 1.520 ;
        RECT  3.770 1.280 4.010 3.370 ;
        RECT  4.010 2.380 4.310 2.660 ;
        RECT  4.310 2.380 4.320 2.650 ;
        RECT  4.320 2.390 4.420 2.650 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 1.780 3.320 2.200 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.040 2.390 1.780 2.650 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.210 2.090 ;
        RECT  0.210 1.830 0.350 2.110 ;
        RECT  0.350 1.830 0.460 2.420 ;
        RECT  0.460 1.870 0.590 2.420 ;
        RECT  0.590 1.870 2.240 2.110 ;
        RECT  2.240 1.870 2.480 2.350 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.800 5.440 ;
        RECT  0.800 3.840 0.810 5.440 ;
        RECT  0.810 3.640 1.210 5.440 ;
        RECT  1.210 3.840 1.220 5.440 ;
        RECT  1.220 4.640 2.140 5.440 ;
        RECT  2.140 3.840 2.150 5.440 ;
        RECT  2.150 3.640 2.550 5.440 ;
        RECT  2.550 3.840 2.560 5.440 ;
        RECT  2.560 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.390 0.400 ;
        RECT  1.390 -0.400 1.790 0.910 ;
        RECT  1.790 -0.400 3.340 0.400 ;
        RECT  3.340 -0.400 3.740 0.560 ;
        RECT  3.740 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.350 3.020 4.750 3.980 ;
        RECT  3.220 3.650 4.350 3.890 ;
        RECT  2.980 2.960 3.220 3.890 ;
        RECT  2.820 2.960 2.980 3.360 ;
        RECT  1.880 3.040 2.820 3.280 ;
        RECT  1.480 2.960 1.880 3.360 ;
        RECT  0.590 3.040 1.480 3.280 ;
        RECT  0.190 2.960 0.590 3.360 ;
    END
END AOI21X2

MACRO AOI21X1
    CLASS CORE ;
    FOREIGN AOI21X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI21XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.570 2.920 2.850 3.900 ;
        RECT  1.390 1.310 2.850 1.550 ;
        RECT  2.850 1.310 2.970 3.900 ;
        RECT  2.970 1.310 3.090 3.210 ;
        RECT  3.090 2.950 3.100 3.210 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.050 1.960 2.180 2.410 ;
        RECT  2.180 1.830 2.440 2.410 ;
        RECT  2.440 1.960 2.460 2.410 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.820 0.550 2.470 ;
        RECT  0.550 2.060 0.690 2.460 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 0.970 3.210 ;
        RECT  0.970 2.390 1.120 3.210 ;
        RECT  1.120 2.390 1.210 3.200 ;
        RECT  1.210 2.390 1.550 2.630 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 4.480 1.390 5.440 ;
        RECT  1.390 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 1.230 ;
        RECT  0.170 -0.400 0.570 1.430 ;
        RECT  0.570 -0.400 0.580 1.230 ;
        RECT  0.580 -0.400 2.310 0.400 ;
        RECT  2.310 -0.400 2.710 0.560 ;
        RECT  2.710 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.810 3.490 2.210 3.890 ;
        RECT  0.570 3.570 1.810 3.810 ;
        RECT  0.170 3.490 0.570 3.890 ;
    END
END AOI21X1

MACRO AOI211XL
    CLASS CORE ;
    FOREIGN AOI211XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.390 0.670 1.770 0.910 ;
        RECT  1.770 0.670 1.780 0.960 ;
        RECT  1.780 0.670 2.020 1.350 ;
        RECT  3.050 2.970 3.500 3.210 ;
        RECT  3.500 2.950 3.510 3.210 ;
        RECT  2.020 1.110 3.510 1.350 ;
        RECT  3.510 1.110 3.750 3.210 ;
        RECT  3.750 2.950 3.760 3.210 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.390 1.670 2.650 ;
        RECT  1.670 2.390 2.440 2.660 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.720 1.590 3.100 2.090 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.380 0.820 2.700 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.270 0.870 1.530 ;
        RECT  0.870 1.270 1.210 1.910 ;
        RECT  1.210 1.670 1.710 1.910 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 4.480 1.390 5.440 ;
        RECT  1.390 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.170 0.400 ;
        RECT  0.170 -0.400 0.570 0.810 ;
        RECT  0.570 -0.400 2.330 0.400 ;
        RECT  2.330 -0.400 2.730 0.560 ;
        RECT  2.730 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  0.170 2.970 2.230 3.210 ;
    END
END AOI211XL

MACRO AOI211X4
    CLASS CORE ;
    FOREIGN AOI211X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI211XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.730 1.260 4.750 2.660 ;
        RECT  4.750 1.260 5.170 3.310 ;
        RECT  5.170 1.260 5.260 1.590 ;
        RECT  5.170 2.890 5.520 3.310 ;
        RECT  5.260 1.190 5.660 1.590 ;
        RECT  5.520 2.900 5.720 3.300 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.390 1.850 2.650 ;
        RECT  1.850 2.370 2.250 2.770 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.530 2.150 2.570 2.550 ;
        RECT  2.570 2.150 2.810 3.750 ;
        RECT  2.810 3.510 2.840 3.750 ;
        RECT  2.810 2.150 2.930 2.550 ;
        RECT  2.840 3.510 3.100 3.770 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.390 0.330 2.650 ;
        RECT  0.330 2.370 0.480 2.650 ;
        RECT  0.480 2.370 0.880 2.770 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.260 1.210 1.920 ;
        RECT  1.210 1.680 1.610 1.920 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.880 5.440 ;
        RECT  0.880 4.360 0.890 5.440 ;
        RECT  0.890 4.160 1.290 5.440 ;
        RECT  1.290 4.360 1.300 5.440 ;
        RECT  1.300 4.640 4.690 5.440 ;
        RECT  4.690 4.320 4.700 5.440 ;
        RECT  4.700 4.120 5.100 5.440 ;
        RECT  5.100 4.320 5.110 5.440 ;
        RECT  5.110 4.640 6.020 5.440 ;
        RECT  6.020 4.480 6.420 5.440 ;
        RECT  6.420 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 0.790 ;
        RECT  0.170 -0.400 0.570 0.990 ;
        RECT  0.570 -0.400 0.580 0.790 ;
        RECT  0.580 -0.400 2.110 0.400 ;
        RECT  2.110 -0.400 2.510 0.560 ;
        RECT  2.510 -0.400 4.480 0.400 ;
        RECT  4.480 -0.400 4.490 0.740 ;
        RECT  4.490 -0.400 4.890 0.940 ;
        RECT  4.890 -0.400 4.900 0.740 ;
        RECT  4.900 -0.400 6.010 0.400 ;
        RECT  6.010 -0.400 6.020 0.950 ;
        RECT  6.020 -0.400 6.420 1.440 ;
        RECT  6.420 -0.400 6.430 0.950 ;
        RECT  6.430 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.000 2.310 6.240 3.840 ;
        RECT  5.810 2.310 6.000 2.550 ;
        RECT  4.320 3.600 6.000 3.840 ;
        RECT  5.410 2.150 5.810 2.550 ;
        RECT  4.080 1.500 4.320 3.840 ;
        RECT  4.050 1.500 4.080 1.740 ;
        RECT  3.900 2.900 4.080 3.300 ;
        RECT  3.810 0.970 4.050 1.740 ;
        RECT  3.500 2.150 3.800 2.550 ;
        RECT  3.290 1.000 3.500 3.150 ;
        RECT  3.260 1.000 3.290 3.230 ;
        RECT  2.990 1.000 3.260 1.400 ;
        RECT  3.050 2.830 3.260 3.230 ;
        RECT  1.770 1.160 2.990 1.400 ;
        RECT  1.610 3.050 2.010 3.550 ;
        RECT  1.530 1.000 1.770 1.400 ;
        RECT  0.570 3.050 1.610 3.290 ;
        RECT  0.170 3.050 0.570 3.550 ;
    END
END AOI211X4

MACRO AOI211X2
    CLASS CORE ;
    FOREIGN AOI211X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI211XL ;
    SIZE 5.940 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  0.170 0.900 0.570 1.300 ;
        RECT  0.570 1.060 2.730 1.300 ;
        RECT  2.730 0.900 3.870 1.300 ;
        RECT  4.030 2.950 4.430 3.380 ;
        RECT  4.430 2.950 4.840 3.210 ;
        RECT  4.840 2.940 5.080 3.210 ;
        RECT  3.870 0.980 5.110 1.220 ;
        RECT  5.080 2.940 5.350 3.200 ;
        RECT  5.110 0.900 5.350 1.300 ;
        RECT  5.350 0.900 5.510 3.200 ;
        RECT  5.510 0.980 5.590 3.200 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.390 3.010 2.650 ;
        RECT  3.010 2.240 3.100 2.650 ;
        RECT  3.100 2.240 3.210 2.640 ;
        RECT  3.210 1.820 3.450 2.640 ;
        RECT  3.450 1.820 4.830 2.060 ;
        RECT  4.830 1.820 5.070 2.230 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.820 2.330 4.500 2.670 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.790 2.400 1.520 2.640 ;
        RECT  1.520 2.390 1.780 2.650 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.460 1.560 0.620 1.950 ;
        RECT  0.620 1.560 0.860 2.080 ;
        RECT  0.860 1.830 1.120 2.090 ;
        RECT  1.120 1.830 2.180 2.080 ;
        RECT  2.180 1.830 2.420 2.910 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.780 5.440 ;
        RECT  0.780 4.130 0.790 5.440 ;
        RECT  0.790 3.930 1.190 5.440 ;
        RECT  1.190 4.130 1.200 5.440 ;
        RECT  1.200 4.640 2.140 5.440 ;
        RECT  2.140 4.130 2.150 5.440 ;
        RECT  2.150 3.930 2.550 5.440 ;
        RECT  2.550 4.130 2.560 5.440 ;
        RECT  2.560 4.640 5.940 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.450 0.400 ;
        RECT  1.450 -0.400 1.850 0.560 ;
        RECT  1.850 -0.400 4.290 0.400 ;
        RECT  4.290 -0.400 4.690 0.560 ;
        RECT  4.690 -0.400 5.940 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  5.250 3.750 5.650 4.150 ;
        RECT  3.290 3.750 5.250 3.990 ;
        RECT  3.050 3.150 3.290 3.990 ;
        RECT  0.170 3.150 3.050 3.390 ;
    END
END AOI211X2

MACRO AOI211X1
    CLASS CORE ;
    FOREIGN AOI211X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AOI211XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  1.390 0.680 1.680 0.920 ;
        RECT  1.680 0.680 1.920 1.160 ;
        RECT  2.910 2.850 3.410 3.830 ;
        RECT  3.410 2.660 3.510 3.830 ;
        RECT  1.920 0.920 3.510 1.160 ;
        RECT  3.510 0.920 3.640 3.830 ;
        RECT  3.640 0.920 3.750 3.780 ;
        RECT  3.750 2.990 3.760 3.780 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 2.370 1.930 2.660 ;
        RECT  1.930 2.290 2.330 2.690 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.630 1.540 3.190 2.100 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 2.040 0.550 2.670 ;
        RECT  0.550 2.260 0.810 2.660 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.270 0.870 1.530 ;
        RECT  0.870 1.270 1.120 1.750 ;
        RECT  1.120 1.510 1.140 1.750 ;
        RECT  1.140 1.510 1.540 1.910 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.920 5.440 ;
        RECT  0.920 3.970 0.930 5.440 ;
        RECT  0.930 3.850 1.330 5.440 ;
        RECT  1.330 3.970 1.340 5.440 ;
        RECT  1.340 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.160 0.400 ;
        RECT  0.160 -0.400 0.170 0.800 ;
        RECT  0.170 -0.400 0.570 0.920 ;
        RECT  0.570 -0.400 0.580 0.800 ;
        RECT  0.580 -0.400 2.210 0.400 ;
        RECT  2.210 -0.400 2.610 0.560 ;
        RECT  2.610 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.690 3.210 2.090 4.190 ;
        RECT  0.570 3.220 1.690 3.460 ;
        RECT  0.170 3.210 0.570 4.190 ;
    END
END AOI211X1

MACRO ANTENNA
    CLASS CORE ;
    FOREIGN ANTENNA 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.320 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.260 0.870 1.880 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.320 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.320 0.400 ;
        END
    END GND
END ANTENNA

MACRO AND4XL
    CLASS CORE ;
    FOREIGN AND4XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.380 0.640 3.480 0.880 ;
        RECT  3.480 0.640 3.720 3.300 ;
        RECT  3.720 0.640 3.760 0.970 ;
        RECT  3.760 0.640 3.780 0.880 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.670 1.770 3.110 2.360 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.150 2.380 1.880 2.760 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 0.920 2.090 ;
        RECT  0.920 1.580 1.400 2.090 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.160 1.180 0.660 1.540 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.840 5.440 ;
        RECT  0.840 4.480 0.920 5.440 ;
        RECT  0.920 4.460 2.340 5.440 ;
        RECT  2.340 4.480 2.990 5.440 ;
        RECT  2.990 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 2.480 0.400 ;
        RECT  2.480 -0.400 2.490 0.660 ;
        RECT  2.490 -0.400 2.890 0.860 ;
        RECT  2.890 -0.400 2.900 0.660 ;
        RECT  2.900 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.390 1.140 3.030 1.380 ;
        RECT  2.240 1.140 2.390 3.330 ;
        RECT  2.240 3.720 2.320 3.960 ;
        RECT  2.150 1.140 2.240 3.960 ;
        RECT  1.920 1.140 2.150 1.380 ;
        RECT  2.000 3.090 2.150 3.960 ;
        RECT  0.850 3.090 2.000 3.330 ;
        RECT  1.920 3.720 2.000 3.960 ;
        RECT  1.680 0.640 1.920 1.380 ;
        RECT  0.180 0.640 1.680 0.880 ;
        RECT  0.450 3.020 0.850 3.330 ;
    END
END AND4XL

MACRO AND4X4
    CLASS CORE ;
    FOREIGN AND4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AND4XL ;
    SIZE 6.600 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.980 1.070 5.380 1.470 ;
        RECT  5.380 1.230 5.390 1.470 ;
        RECT  5.390 1.230 5.630 4.360 ;
        RECT  5.630 2.940 5.830 4.340 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  3.940 2.290 4.510 2.940 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.840 2.390 2.860 2.650 ;
        RECT  2.860 2.390 3.100 2.900 ;
        RECT  3.100 2.660 3.230 2.900 ;
        RECT  3.230 2.660 3.630 3.060 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.180 1.830 2.240 2.090 ;
        RECT  2.240 1.830 2.440 3.010 ;
        RECT  2.440 1.840 2.480 3.010 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 1.120 2.650 ;
        RECT  1.120 2.390 1.450 2.630 ;
        RECT  1.450 2.170 1.720 2.630 ;
        RECT  1.720 2.170 1.850 2.570 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.230 5.440 ;
        RECT  1.230 3.900 1.240 5.440 ;
        RECT  1.240 3.410 1.640 5.440 ;
        RECT  1.640 3.900 1.650 5.440 ;
        RECT  1.650 4.640 2.810 5.440 ;
        RECT  2.810 4.010 2.820 5.440 ;
        RECT  2.820 3.890 3.220 5.440 ;
        RECT  3.220 4.010 3.230 5.440 ;
        RECT  3.230 4.640 4.500 5.440 ;
        RECT  4.500 4.010 4.510 5.440 ;
        RECT  4.510 3.890 4.910 5.440 ;
        RECT  4.910 4.010 4.920 5.440 ;
        RECT  4.920 4.640 6.110 5.440 ;
        RECT  6.110 2.940 6.350 5.440 ;
        RECT  6.350 4.640 6.600 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 3.680 0.400 ;
        RECT  3.680 -0.400 3.690 0.990 ;
        RECT  3.690 -0.400 4.660 1.480 ;
        RECT  4.660 -0.400 4.670 0.990 ;
        RECT  4.670 -0.400 5.900 0.400 ;
        RECT  5.900 -0.400 5.910 1.330 ;
        RECT  5.910 -0.400 6.310 1.530 ;
        RECT  6.310 -0.400 6.320 1.330 ;
        RECT  6.320 -0.400 6.600 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  4.780 1.750 5.020 3.610 ;
        RECT  3.090 1.750 4.780 1.990 ;
        RECT  4.110 3.370 4.780 3.610 ;
        RECT  3.710 3.360 4.110 4.340 ;
        RECT  2.360 3.370 3.710 3.610 ;
        RECT  2.850 1.220 3.090 1.990 ;
        RECT  1.990 1.220 2.850 1.460 ;
        RECT  1.960 3.300 2.360 4.280 ;
        RECT  1.590 1.060 1.990 1.460 ;
    END
END AND4X4

MACRO AND4X2
    CLASS CORE ;
    FOREIGN AND4X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AND4XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.200 1.100 3.520 1.530 ;
        RECT  3.520 1.100 3.600 1.540 ;
        RECT  3.600 1.270 3.760 1.540 ;
        RECT  3.760 1.300 4.050 1.540 ;
        RECT  4.050 1.300 4.290 3.800 ;
        RECT  4.290 2.640 4.450 3.800 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.390 2.380 2.400 2.660 ;
        RECT  2.400 2.380 2.800 2.840 ;
        RECT  2.800 2.380 3.190 2.660 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.830 1.530 2.090 ;
        RECT  1.530 1.830 1.780 2.450 ;
        RECT  1.780 2.050 2.010 2.450 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.950 0.870 3.210 ;
        RECT  0.870 2.290 1.110 3.210 ;
        RECT  1.110 2.950 1.120 3.210 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.460 0.460 2.090 ;
        RECT  0.460 1.460 0.500 1.880 ;
        RECT  0.500 1.470 0.810 1.870 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.170 5.440 ;
        RECT  0.170 4.480 1.790 5.440 ;
        RECT  1.790 4.640 3.230 5.440 ;
        RECT  3.230 4.480 3.630 5.440 ;
        RECT  3.630 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 2.370 0.400 ;
        RECT  2.370 -0.400 2.770 0.560 ;
        RECT  2.770 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.530 1.810 3.770 3.600 ;
        RECT  2.530 1.810 3.530 2.050 ;
        RECT  2.600 3.360 3.530 3.600 ;
        RECT  2.200 3.360 2.600 3.760 ;
        RECT  2.290 0.860 2.530 2.050 ;
        RECT  1.400 0.860 2.290 1.100 ;
        RECT  1.180 3.490 2.200 3.730 ;
        RECT  1.160 0.670 1.400 1.100 ;
        RECT  0.780 3.490 1.180 3.890 ;
        RECT  0.170 0.670 1.160 0.910 ;
    END
END AND4X2

MACRO AND4X1
    CLASS CORE ;
    FOREIGN AND4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AND4XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.400 2.940 3.480 3.340 ;
        RECT  3.320 0.670 3.480 0.910 ;
        RECT  3.480 0.670 3.720 3.340 ;
        RECT  3.720 0.670 3.750 0.970 ;
        RECT  3.750 0.710 3.760 0.970 ;
        RECT  3.720 2.940 3.800 3.340 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.760 1.830 3.110 2.480 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.310 2.360 1.980 2.800 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 1.830 0.920 2.090 ;
        RECT  0.920 1.630 1.400 2.100 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.160 1.180 0.660 1.540 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.840 5.440 ;
        RECT  0.840 4.480 0.920 5.440 ;
        RECT  0.920 4.460 2.340 5.440 ;
        RECT  2.340 4.480 2.990 5.440 ;
        RECT  2.990 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 2.490 0.400 ;
        RECT  2.490 -0.400 2.890 0.560 ;
        RECT  2.890 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.490 1.280 3.030 1.520 ;
        RECT  2.320 1.280 2.490 3.340 ;
        RECT  2.250 1.280 2.320 4.040 ;
        RECT  1.920 1.280 2.250 1.520 ;
        RECT  1.920 3.100 2.250 4.040 ;
        RECT  1.680 0.680 1.920 1.520 ;
        RECT  0.850 3.100 1.920 3.340 ;
        RECT  0.180 0.680 1.680 0.920 ;
        RECT  0.450 2.940 0.850 3.340 ;
    END
END AND4X1

MACRO AND3XL
    CLASS CORE ;
    FOREIGN AND3XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.660 3.740 2.890 4.110 ;
        RECT  2.750 1.270 2.890 1.870 ;
        RECT  2.890 1.270 3.130 4.110 ;
        RECT  3.130 1.270 3.140 1.870 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.370 1.850 1.520 2.430 ;
        RECT  1.520 1.830 1.610 2.430 ;
        RECT  1.610 1.830 1.780 2.090 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.810 2.740 1.210 3.220 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.160 3.510 0.800 3.800 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.800 5.440 ;
        RECT  1.800 4.480 2.030 5.440 ;
        RECT  2.030 3.260 2.270 5.440 ;
        RECT  2.270 3.260 2.370 3.500 ;
        RECT  2.370 2.970 2.610 3.500 ;
        RECT  2.270 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.970 0.400 ;
        RECT  1.970 -0.400 2.370 0.560 ;
        RECT  2.370 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.180 1.190 2.420 2.690 ;
        RECT  1.140 1.190 2.180 1.430 ;
        RECT  2.090 2.450 2.180 2.690 ;
        RECT  1.850 2.450 2.090 2.950 ;
        RECT  1.730 2.710 1.850 2.950 ;
        RECT  1.520 2.710 1.730 3.730 ;
        RECT  1.490 2.710 1.520 4.360 ;
        RECT  1.280 3.490 1.490 4.360 ;
        RECT  0.170 4.120 1.280 4.360 ;
        RECT  0.900 0.640 1.140 1.430 ;
        RECT  0.170 0.640 0.900 0.880 ;
    END
END AND3XL

MACRO AND3X4
    CLASS CORE ;
    FOREIGN AND3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AND3XL ;
    SIZE 5.280 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  4.030 0.730 4.070 1.710 ;
        RECT  4.030 2.920 4.080 4.180 ;
        RECT  4.070 0.730 4.080 2.660 ;
        RECT  4.080 0.730 4.270 4.180 ;
        RECT  4.270 0.730 4.430 4.160 ;
        RECT  4.430 0.730 4.510 2.660 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.750 2.250 3.190 2.660 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  2.040 2.620 2.120 3.020 ;
        RECT  2.120 2.620 2.180 3.200 ;
        RECT  2.180 2.620 2.440 3.210 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.380 1.320 2.660 ;
        RECT  1.320 2.040 1.720 2.660 ;
        RECT  1.720 2.380 1.730 2.660 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.660 5.440 ;
        RECT  1.660 4.210 1.670 5.440 ;
        RECT  1.670 4.010 2.070 5.440 ;
        RECT  2.070 4.210 2.080 5.440 ;
        RECT  2.080 4.640 3.180 5.440 ;
        RECT  3.180 4.210 3.190 5.440 ;
        RECT  3.190 4.010 3.590 5.440 ;
        RECT  3.590 4.210 3.600 5.440 ;
        RECT  3.600 4.640 4.700 5.440 ;
        RECT  4.700 3.700 4.710 5.440 ;
        RECT  4.710 3.210 5.110 5.440 ;
        RECT  5.110 3.700 5.120 5.440 ;
        RECT  5.120 4.640 5.280 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 3.100 0.400 ;
        RECT  3.100 -0.400 3.110 0.830 ;
        RECT  3.110 -0.400 3.510 1.030 ;
        RECT  3.510 -0.400 3.520 0.830 ;
        RECT  3.520 -0.400 4.790 0.400 ;
        RECT  4.790 -0.400 5.030 1.710 ;
        RECT  5.030 -0.400 5.280 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  3.700 2.150 3.800 2.630 ;
        RECT  3.460 1.310 3.700 3.730 ;
        RECT  2.730 1.310 3.460 1.550 ;
        RECT  2.830 3.490 3.460 3.730 ;
        RECT  2.430 3.490 2.830 3.890 ;
        RECT  2.490 1.220 2.730 1.550 ;
        RECT  1.740 1.220 2.490 1.460 ;
        RECT  1.300 3.490 2.430 3.730 ;
        RECT  1.340 1.060 1.740 1.460 ;
        RECT  0.900 3.490 1.300 3.890 ;
    END
END AND3X4

MACRO AND3X2
    CLASS CORE ;
    FOREIGN AND3X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AND3XL ;
    SIZE 3.960 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.390 3.190 3.500 4.170 ;
        RECT  3.500 2.950 3.510 4.170 ;
        RECT  3.390 1.110 3.510 1.510 ;
        RECT  3.510 1.110 3.750 4.170 ;
        RECT  3.750 2.950 3.760 4.170 ;
        RECT  3.760 3.190 3.790 4.170 ;
        RECT  3.750 1.110 3.790 1.510 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.520 1.820 1.930 2.100 ;
        RECT  1.930 1.670 2.330 2.100 ;
        RECT  2.330 1.820 2.340 2.100 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 1.560 2.800 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.820 0.530 2.090 ;
        RECT  0.530 1.660 0.930 2.090 ;
        RECT  0.930 1.820 0.940 2.090 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.930 5.440 ;
        RECT  0.930 4.480 1.330 5.440 ;
        RECT  1.330 4.640 2.570 5.440 ;
        RECT  2.570 4.480 2.970 5.440 ;
        RECT  2.970 4.640 3.960 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 2.570 0.400 ;
        RECT  2.570 -0.400 2.970 0.560 ;
        RECT  2.970 -0.400 3.960 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.950 1.810 3.110 2.210 ;
        RECT  2.710 1.070 2.950 3.360 ;
        RECT  1.190 1.070 2.710 1.310 ;
        RECT  2.090 3.120 2.710 3.360 ;
        RECT  1.690 3.120 2.090 3.730 ;
        RECT  0.170 3.490 1.690 3.730 ;
        RECT  0.950 0.890 1.190 1.310 ;
        RECT  0.270 0.890 0.950 1.130 ;
    END
END AND3X2

MACRO AND3X1
    CLASS CORE ;
    FOREIGN AND3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AND3XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.770 3.970 2.850 4.370 ;
        RECT  2.760 1.270 2.850 1.820 ;
        RECT  2.840 0.710 2.850 0.970 ;
        RECT  2.850 0.710 3.010 4.370 ;
        RECT  3.010 0.710 3.090 4.210 ;
        RECT  3.090 0.710 3.100 0.970 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.320 1.840 1.520 2.440 ;
        RECT  1.520 1.830 1.560 2.440 ;
        RECT  1.560 1.830 1.780 2.090 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.810 2.710 1.210 3.220 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 3.510 0.760 3.850 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.840 5.440 ;
        RECT  1.840 4.480 2.000 5.440 ;
        RECT  2.000 3.450 2.240 5.440 ;
        RECT  2.240 3.450 2.360 3.690 ;
        RECT  2.360 2.890 2.600 3.690 ;
        RECT  2.240 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 2.020 0.400 ;
        RECT  2.020 -0.400 2.420 0.560 ;
        RECT  2.420 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.190 1.310 2.430 2.610 ;
        RECT  1.060 1.310 2.190 1.550 ;
        RECT  2.080 2.370 2.190 2.610 ;
        RECT  1.840 2.370 2.080 3.010 ;
        RECT  1.720 2.770 1.840 3.010 ;
        RECT  1.560 2.770 1.720 4.170 ;
        RECT  1.480 2.770 1.560 4.370 ;
        RECT  1.320 3.930 1.480 4.370 ;
        RECT  0.170 4.130 1.320 4.370 ;
        RECT  0.820 0.640 1.060 1.550 ;
        RECT  0.170 0.640 0.820 0.880 ;
    END
END AND3X1

MACRO AND2XL
    CLASS CORE ;
    FOREIGN AND2XL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.150 1.250 2.390 3.520 ;
        RECT  2.390 2.390 2.440 2.650 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.380 1.250 2.950 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.810 0.510 2.450 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.390 5.440 ;
        RECT  0.390 4.480 1.370 5.440 ;
        RECT  1.370 4.640 2.640 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.360 0.400 ;
        RECT  1.360 -0.400 1.760 0.560 ;
        RECT  1.760 -0.400 2.640 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.580 0.860 1.820 3.480 ;
        RECT  1.080 0.860 1.580 1.100 ;
        RECT  0.450 3.240 1.580 3.480 ;
        RECT  0.840 0.670 1.080 1.100 ;
        RECT  0.180 0.670 0.840 0.910 ;
    END
END AND2XL

MACRO AND2X4
    CLASS CORE ;
    FOREIGN AND2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AND2XL ;
    SIZE 4.620 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.500 2.870 2.750 3.830 ;
        RECT  2.750 2.380 2.790 3.830 ;
        RECT  2.530 1.150 2.790 1.550 ;
        RECT  2.790 1.150 2.900 3.830 ;
        RECT  2.900 1.150 3.030 3.780 ;
        RECT  3.030 2.380 3.190 3.780 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.940 1.120 3.210 ;
        RECT  1.120 2.940 1.420 3.200 ;
        RECT  1.420 2.220 1.660 3.200 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 1.030 2.110 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.240 5.440 ;
        RECT  0.240 3.770 0.250 5.440 ;
        RECT  0.250 3.570 0.650 5.440 ;
        RECT  0.650 3.770 0.660 5.440 ;
        RECT  0.660 4.640 1.800 5.440 ;
        RECT  1.800 4.480 2.200 5.440 ;
        RECT  2.200 4.640 3.140 5.440 ;
        RECT  3.140 4.340 3.150 5.440 ;
        RECT  3.150 4.140 3.550 5.440 ;
        RECT  3.550 4.340 3.560 5.440 ;
        RECT  3.560 4.640 4.620 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.850 0.400 ;
        RECT  1.850 -0.400 1.860 0.670 ;
        RECT  1.860 -0.400 2.260 0.870 ;
        RECT  2.260 -0.400 2.270 0.670 ;
        RECT  2.270 -0.400 3.140 0.400 ;
        RECT  3.140 -0.400 3.150 0.670 ;
        RECT  3.150 -0.400 3.550 0.870 ;
        RECT  3.550 -0.400 3.560 0.670 ;
        RECT  3.560 -0.400 4.620 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  2.180 1.860 2.510 2.100 ;
        RECT  1.940 1.150 2.180 3.810 ;
        RECT  1.040 1.150 1.940 1.390 ;
        RECT  1.390 3.570 1.940 3.810 ;
        RECT  0.990 3.490 1.390 3.890 ;
        RECT  0.640 0.990 1.040 1.390 ;
    END
END AND2X4

MACRO AND2X2
    CLASS CORE ;
    FOREIGN AND2X2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AND2XL ;
    SIZE 3.300 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.680 1.150 2.690 3.450 ;
        RECT  2.690 0.660 3.090 3.940 ;
        RECT  3.090 0.820 3.100 3.940 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.290 3.520 1.520 4.110 ;
        RECT  1.520 3.510 1.690 4.110 ;
        RECT  1.690 3.510 1.780 3.770 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.820 0.550 2.450 ;
        RECT  0.550 1.830 0.850 2.230 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.160 5.440 ;
        RECT  0.160 3.690 0.170 5.440 ;
        RECT  0.170 3.490 0.570 5.440 ;
        RECT  0.570 3.690 0.580 5.440 ;
        RECT  0.580 4.640 1.870 5.440 ;
        RECT  1.870 4.480 2.270 5.440 ;
        RECT  2.270 4.640 3.300 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.920 0.400 ;
        RECT  1.920 -0.400 1.930 0.970 ;
        RECT  1.930 -0.400 2.330 1.460 ;
        RECT  2.330 -0.400 2.340 0.970 ;
        RECT  2.340 -0.400 3.300 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.370 1.840 2.410 2.240 ;
        RECT  1.370 2.830 1.450 3.230 ;
        RECT  1.130 1.120 1.370 3.230 ;
        RECT  0.980 1.120 1.130 1.360 ;
        RECT  1.050 2.830 1.130 3.230 ;
        RECT  0.580 0.960 0.980 1.360 ;
    END
END AND2X2

MACRO AND2X1
    CLASS CORE ;
    FOREIGN AND2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ AND2XL ;
    SIZE 2.640 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  2.140 1.200 2.380 3.520 ;
        RECT  2.380 2.390 2.440 2.650 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.830 2.390 1.220 2.960 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.160 1.810 0.520 2.460 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.490 5.440 ;
        RECT  0.490 4.480 1.470 5.440 ;
        RECT  1.470 4.640 2.640 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.360 0.400 ;
        RECT  1.360 -0.400 1.760 0.560 ;
        RECT  1.760 -0.400 2.640 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  1.590 0.860 1.830 3.480 ;
        RECT  1.070 0.860 1.590 1.100 ;
        RECT  0.450 3.240 1.590 3.480 ;
        RECT  0.830 0.670 1.070 1.100 ;
        RECT  0.180 0.670 0.830 0.910 ;
    END
END AND2X1

MACRO ADDHXL
    CLASS CORE ;
    FOREIGN ADDHXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.920 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 2.950 3.510 3.220 ;
        RECT  3.510 2.950 3.750 3.520 ;
        RECT  3.570 1.190 3.810 1.860 ;
        RECT  3.750 2.950 4.470 3.220 ;
        RECT  3.810 1.620 4.470 1.860 ;
        RECT  4.470 1.620 4.710 3.220 ;
        RECT  4.710 2.950 4.720 3.220 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  7.240 1.390 7.370 1.790 ;
        RECT  7.370 1.390 7.460 1.830 ;
        RECT  7.350 2.980 7.470 3.380 ;
        RECT  7.460 1.390 7.470 2.090 ;
        RECT  7.470 1.390 7.640 3.380 ;
        RECT  7.640 1.550 7.710 3.380 ;
        RECT  7.710 1.830 7.720 2.090 ;
        RECT  7.710 2.980 7.750 3.380 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.840 2.430 2.750 2.830 ;
        RECT  2.750 2.430 2.990 3.210 ;
        RECT  2.990 2.430 3.230 4.290 ;
        RECT  3.230 2.430 3.570 2.670 ;
        RECT  3.570 2.140 3.810 2.670 ;
        RECT  3.810 2.140 4.190 2.380 ;
        RECT  3.230 4.050 5.510 4.290 ;
        RECT  5.510 3.820 5.750 4.290 ;
        RECT  5.750 3.820 6.120 4.060 ;
        RECT  6.120 3.660 6.520 4.060 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  5.500 1.820 5.510 2.100 ;
        RECT  5.510 1.820 5.750 2.590 ;
        RECT  5.750 1.820 6.400 2.100 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.980 5.440 ;
        RECT  0.980 4.480 1.380 5.440 ;
        RECT  1.380 4.640 6.020 5.440 ;
        RECT  6.020 4.480 7.000 5.440 ;
        RECT  7.000 4.640 7.920 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.050 0.400 ;
        RECT  1.050 -0.400 1.450 0.560 ;
        RECT  1.450 -0.400 5.080 0.400 ;
        RECT  5.080 -0.400 5.480 0.560 ;
        RECT  5.480 -0.400 7.170 0.400 ;
        RECT  7.170 -0.400 7.570 0.560 ;
        RECT  7.570 -0.400 7.920 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  6.760 1.280 7.000 3.210 ;
        RECT  6.330 1.280 6.760 1.520 ;
        RECT  6.220 2.970 6.760 3.210 ;
        RECT  5.820 2.970 6.220 3.370 ;
        RECT  4.990 1.100 5.230 3.770 ;
        RECT  4.330 1.100 4.990 1.340 ;
        RECT  4.190 3.530 4.990 3.770 ;
        RECT  4.090 0.670 4.330 1.340 ;
        RECT  3.290 0.670 4.090 0.910 ;
        RECT  3.050 0.670 3.290 2.140 ;
        RECT  1.440 1.900 3.050 2.140 ;
        RECT  2.530 0.700 2.770 1.100 ;
        RECT  2.470 3.490 2.710 4.180 ;
        RECT  0.920 1.380 2.680 1.620 ;
        RECT  0.400 0.860 2.530 1.100 ;
        RECT  0.570 3.940 2.470 4.180 ;
        RECT  1.540 3.380 2.050 3.620 ;
        RECT  1.300 2.980 1.540 3.620 ;
        RECT  1.200 1.900 1.440 2.700 ;
        RECT  0.920 2.980 1.300 3.220 ;
        RECT  0.680 1.380 0.920 3.220 ;
        RECT  0.400 3.500 0.570 4.180 ;
        RECT  0.160 0.860 0.400 4.180 ;
    END
END ADDHXL

MACRO ADDHX4
    CLASS CORE ;
    FOREIGN ADDHX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ ADDHXL ;
    SIZE 20.460 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  5.570 2.730 6.710 3.150 ;
        RECT  6.360 1.240 6.710 1.660 ;
        RECT  6.710 1.240 6.810 3.150 ;
        RECT  6.810 1.240 6.990 3.170 ;
        RECT  6.990 1.250 7.050 3.170 ;
        RECT  7.050 1.250 7.130 3.330 ;
        RECT  7.130 1.250 7.150 2.660 ;
        RECT  7.150 1.250 8.030 1.650 ;
        RECT  8.030 1.240 9.070 1.660 ;
        RECT  9.070 0.640 9.270 1.660 ;
        RECT  9.270 0.640 9.420 1.620 ;
        RECT  7.130 2.930 11.940 3.330 ;
        RECT  9.420 0.640 12.100 0.980 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  19.220 2.380 19.250 3.760 ;
        RECT  19.250 2.380 19.690 3.780 ;
        RECT  19.690 2.380 19.880 2.780 ;
        RECT  18.600 1.190 19.880 1.590 ;
        RECT  19.880 1.190 20.280 2.780 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.410 2.350 9.440 2.590 ;
        RECT  9.440 2.350 9.540 2.650 ;
        RECT  9.540 1.890 9.700 2.650 ;
        RECT  9.700 1.890 9.780 2.640 ;
        RECT  9.780 1.890 12.090 2.130 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  13.790 1.990 14.060 2.230 ;
        RECT  14.060 1.830 14.320 2.230 ;
        RECT  14.320 1.990 17.910 2.230 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.300 5.440 ;
        RECT  0.300 3.590 0.310 5.440 ;
        RECT  0.310 2.840 0.710 5.440 ;
        RECT  0.710 3.590 0.720 5.440 ;
        RECT  0.720 4.640 1.840 5.440 ;
        RECT  1.840 3.740 1.850 5.440 ;
        RECT  1.850 3.260 2.250 5.440 ;
        RECT  2.250 3.740 2.260 5.440 ;
        RECT  2.260 4.640 3.390 5.440 ;
        RECT  3.390 4.480 3.790 5.440 ;
        RECT  3.790 4.640 4.860 5.440 ;
        RECT  4.860 4.480 5.260 5.440 ;
        RECT  5.260 4.640 12.180 5.440 ;
        RECT  12.180 4.480 12.580 5.440 ;
        RECT  12.580 4.640 13.770 5.440 ;
        RECT  13.770 4.480 14.170 5.440 ;
        RECT  14.170 4.640 15.320 5.440 ;
        RECT  15.320 3.810 15.330 5.440 ;
        RECT  15.330 3.610 15.730 5.440 ;
        RECT  15.730 3.810 15.740 5.440 ;
        RECT  15.740 4.640 16.860 5.440 ;
        RECT  16.860 3.810 16.870 5.440 ;
        RECT  16.870 3.610 17.270 5.440 ;
        RECT  17.270 3.810 17.280 5.440 ;
        RECT  17.280 4.640 18.510 5.440 ;
        RECT  18.510 4.030 18.910 5.440 ;
        RECT  18.910 4.640 19.900 5.440 ;
        RECT  19.900 4.030 20.300 5.440 ;
        RECT  20.300 4.640 20.460 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.980 0.400 ;
        RECT  0.980 -0.400 0.990 0.900 ;
        RECT  0.990 -0.400 1.390 1.100 ;
        RECT  1.390 -0.400 1.400 0.900 ;
        RECT  1.400 -0.400 2.270 0.400 ;
        RECT  2.270 -0.400 2.280 0.900 ;
        RECT  2.280 -0.400 2.680 1.100 ;
        RECT  2.680 -0.400 2.690 0.900 ;
        RECT  2.690 -0.400 3.650 0.400 ;
        RECT  3.650 -0.400 4.050 0.560 ;
        RECT  4.050 -0.400 5.170 0.400 ;
        RECT  5.170 -0.400 5.570 0.560 ;
        RECT  5.570 -0.400 14.030 0.400 ;
        RECT  14.030 -0.400 14.040 0.830 ;
        RECT  14.040 -0.400 14.440 0.950 ;
        RECT  14.440 -0.400 14.450 0.830 ;
        RECT  14.450 -0.400 15.340 0.400 ;
        RECT  15.340 -0.400 15.350 0.830 ;
        RECT  15.350 -0.400 15.750 1.030 ;
        RECT  15.750 -0.400 15.760 0.830 ;
        RECT  15.760 -0.400 16.680 0.400 ;
        RECT  16.680 -0.400 16.690 0.830 ;
        RECT  16.690 -0.400 17.090 1.030 ;
        RECT  17.090 -0.400 17.100 0.830 ;
        RECT  17.100 -0.400 17.970 0.400 ;
        RECT  17.970 -0.400 17.980 0.710 ;
        RECT  17.980 -0.400 18.380 0.910 ;
        RECT  18.380 -0.400 18.390 0.710 ;
        RECT  18.390 -0.400 19.230 0.400 ;
        RECT  19.230 -0.400 19.240 0.710 ;
        RECT  19.240 -0.400 19.640 0.910 ;
        RECT  19.640 -0.400 19.650 0.710 ;
        RECT  19.650 -0.400 20.460 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  18.820 1.870 19.640 2.110 ;
        RECT  18.580 1.870 18.820 2.750 ;
        RECT  13.370 2.510 18.580 2.750 ;
        RECT  17.640 3.020 18.040 3.980 ;
        RECT  17.310 1.310 17.710 1.710 ;
        RECT  16.500 3.030 17.640 3.270 ;
        RECT  16.420 1.390 17.310 1.630 ;
        RECT  16.100 3.020 16.500 3.980 ;
        RECT  16.020 1.310 16.420 1.710 ;
        RECT  14.960 3.030 16.100 3.270 ;
        RECT  15.080 1.390 16.020 1.630 ;
        RECT  14.680 1.310 15.080 1.710 ;
        RECT  14.560 3.020 14.960 3.980 ;
        RECT  13.770 1.310 14.680 1.550 ;
        RECT  13.910 3.030 14.560 3.270 ;
        RECT  13.670 3.030 13.910 3.850 ;
        RECT  13.530 0.690 13.770 1.550 ;
        RECT  12.620 3.610 13.670 3.850 ;
        RECT  12.620 0.690 13.530 0.930 ;
        RECT  13.160 2.510 13.370 3.210 ;
        RECT  12.970 1.300 13.160 3.210 ;
        RECT  12.920 1.300 12.970 2.750 ;
        RECT  12.380 0.690 12.620 3.850 ;
        RECT  9.770 1.330 12.380 1.570 ;
        RECT  11.300 3.610 12.380 3.850 ;
        RECT  10.900 3.610 11.300 4.110 ;
        RECT  9.870 3.610 10.900 3.850 ;
        RECT  9.760 3.610 9.870 4.030 ;
        RECT  9.360 3.610 9.760 4.110 ;
        RECT  6.390 3.610 9.360 3.850 ;
        RECT  6.090 0.650 8.730 0.890 ;
        RECT  5.760 4.130 8.220 4.370 ;
        RECT  6.150 3.420 6.390 3.850 ;
        RECT  3.630 3.420 6.150 3.660 ;
        RECT  5.850 0.650 6.090 1.120 ;
        RECT  5.970 1.670 6.090 2.070 ;
        RECT  4.840 1.660 5.970 2.080 ;
        RECT  3.350 0.880 5.850 1.120 ;
        RECT  5.520 3.940 5.760 4.370 ;
        RECT  3.000 3.940 5.520 4.180 ;
        RECT  4.570 1.380 4.840 2.080 ;
        RECT  4.560 1.380 4.570 3.020 ;
        RECT  4.440 1.380 4.560 3.140 ;
        RECT  4.160 1.660 4.440 3.140 ;
        RECT  4.150 1.660 4.160 3.020 ;
        RECT  3.390 2.230 3.630 3.660 ;
        RECT  3.300 2.230 3.390 2.470 ;
        RECT  3.110 0.880 3.350 1.780 ;
        RECT  1.760 2.070 3.300 2.470 ;
        RECT  2.950 1.380 3.110 1.780 ;
        RECT  3.000 2.740 3.020 3.700 ;
        RECT  2.760 2.740 3.000 4.180 ;
        RECT  2.010 1.540 2.950 1.780 ;
        RECT  2.620 2.740 2.760 3.700 ;
        RECT  1.480 2.750 2.620 2.990 ;
        RECT  1.610 1.380 2.010 1.780 ;
        RECT  1.400 1.540 1.610 1.780 ;
        RECT  1.400 2.740 1.480 3.700 ;
        RECT  1.160 1.540 1.400 3.700 ;
        RECT  1.080 2.740 1.160 3.700 ;
    END
END ADDHX4

MACRO ADDHX2
    CLASS CORE ;
    FOREIGN ADDHX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ ADDHXL ;
    SIZE 13.200 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.410 2.900 3.620 3.140 ;
        RECT  3.620 1.350 3.860 3.140 ;
        RECT  3.860 2.900 4.160 3.140 ;
        RECT  4.160 2.900 4.420 3.210 ;
        RECT  4.420 2.900 4.960 3.140 ;
        RECT  4.960 2.900 5.200 3.870 ;
        RECT  5.200 2.930 5.390 3.220 ;
        RECT  5.390 2.930 5.490 3.200 ;
        RECT  5.490 2.930 6.290 3.170 ;
        RECT  6.290 2.930 6.690 3.330 ;
        RECT  3.860 1.350 6.690 1.590 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.030 1.210 12.090 1.610 ;
        RECT  12.080 2.950 12.130 3.210 ;
        RECT  12.090 1.210 12.130 1.840 ;
        RECT  12.130 1.210 12.370 3.210 ;
        RECT  12.370 1.210 12.430 1.970 ;
        RECT  12.370 2.520 12.670 3.210 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.140 2.350 5.480 2.590 ;
        RECT  5.480 2.350 5.520 2.650 ;
        RECT  5.520 1.930 5.740 2.650 ;
        RECT  5.740 1.930 5.830 2.590 ;
        RECT  5.830 1.930 6.500 2.170 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  8.120 1.830 8.130 2.090 ;
        RECT  8.130 1.830 8.380 2.190 ;
        RECT  8.380 1.950 10.240 2.190 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.300 5.440 ;
        RECT  0.300 4.210 0.310 5.440 ;
        RECT  0.310 4.010 0.710 5.440 ;
        RECT  0.710 4.210 0.720 5.440 ;
        RECT  0.720 4.640 1.830 5.440 ;
        RECT  1.830 4.480 2.230 5.440 ;
        RECT  2.230 4.640 7.150 5.440 ;
        RECT  7.150 4.480 7.550 5.440 ;
        RECT  7.550 4.640 8.780 5.440 ;
        RECT  8.780 4.120 8.790 5.440 ;
        RECT  8.790 3.920 9.190 5.440 ;
        RECT  9.190 4.120 9.200 5.440 ;
        RECT  9.200 4.640 10.260 5.440 ;
        RECT  10.260 4.120 10.270 5.440 ;
        RECT  10.270 3.920 10.670 5.440 ;
        RECT  10.670 4.120 10.680 5.440 ;
        RECT  10.680 4.640 11.650 5.440 ;
        RECT  11.650 4.120 11.660 5.440 ;
        RECT  11.660 3.920 12.060 5.440 ;
        RECT  12.060 4.120 12.070 5.440 ;
        RECT  12.070 4.640 13.200 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.540 0.400 ;
        RECT  0.540 -0.400 0.550 0.910 ;
        RECT  0.550 -0.400 0.950 1.110 ;
        RECT  0.950 -0.400 0.960 0.910 ;
        RECT  0.960 -0.400 1.890 0.400 ;
        RECT  1.890 -0.400 2.290 0.560 ;
        RECT  2.290 -0.400 8.680 0.400 ;
        RECT  8.680 -0.400 8.690 0.790 ;
        RECT  8.690 -0.400 9.090 0.990 ;
        RECT  9.090 -0.400 9.100 0.790 ;
        RECT  9.100 -0.400 9.960 0.400 ;
        RECT  9.960 -0.400 9.970 0.790 ;
        RECT  9.970 -0.400 10.370 0.990 ;
        RECT  10.370 -0.400 10.380 0.790 ;
        RECT  10.380 -0.400 11.410 0.400 ;
        RECT  11.410 -0.400 11.420 0.730 ;
        RECT  11.420 -0.400 11.820 0.930 ;
        RECT  11.820 -0.400 11.830 0.730 ;
        RECT  11.830 -0.400 13.200 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  11.440 2.130 11.840 2.530 ;
        RECT  10.770 2.290 11.440 2.530 ;
        RECT  9.930 2.990 11.320 3.230 ;
        RECT  10.680 1.270 11.080 1.670 ;
        RECT  10.530 2.290 10.770 2.710 ;
        RECT  9.730 1.270 10.680 1.510 ;
        RECT  8.370 2.470 10.530 2.710 ;
        RECT  9.530 2.980 9.930 3.940 ;
        RECT  9.330 1.270 9.730 1.670 ;
        RECT  7.270 3.400 9.530 3.640 ;
        RECT  8.350 1.270 9.330 1.510 ;
        RECT  7.970 2.470 8.370 3.120 ;
        RECT  8.110 0.680 8.350 1.510 ;
        RECT  7.210 0.680 8.110 0.920 ;
        RECT  7.730 2.470 7.970 2.710 ;
        RECT  7.490 1.200 7.730 2.710 ;
        RECT  7.210 3.400 7.270 3.850 ;
        RECT  6.970 0.680 7.210 3.850 ;
        RECT  6.050 0.680 6.970 0.920 ;
        RECT  6.050 3.610 6.970 3.850 ;
        RECT  5.650 0.670 6.050 0.920 ;
        RECT  5.860 3.610 6.050 4.200 ;
        RECT  5.620 3.610 5.860 4.370 ;
        RECT  2.750 4.130 5.620 4.370 ;
        RECT  4.480 0.670 4.700 0.910 ;
        RECT  3.410 3.610 4.540 3.850 ;
        RECT  4.240 0.670 4.480 0.990 ;
        RECT  2.810 0.750 4.240 0.990 ;
        RECT  3.170 3.420 3.410 3.850 ;
        RECT  3.120 1.880 3.350 2.280 ;
        RECT  1.950 3.420 3.170 3.660 ;
        RECT  3.110 1.870 3.120 2.290 ;
        RECT  3.030 1.390 3.110 2.290 ;
        RECT  3.030 2.900 3.050 3.140 ;
        RECT  2.790 1.390 3.030 3.140 ;
        RECT  2.570 0.750 2.810 1.100 ;
        RECT  2.710 1.390 2.790 1.630 ;
        RECT  2.650 2.900 2.790 3.140 ;
        RECT  2.510 3.940 2.750 4.370 ;
        RECT  1.950 0.860 2.570 1.100 ;
        RECT  1.230 3.940 2.510 4.180 ;
        RECT  1.710 0.860 1.950 3.660 ;
        RECT  1.190 1.390 1.710 1.790 ;
        RECT  1.030 2.770 1.710 3.170 ;
        RECT  1.030 2.090 1.430 2.490 ;
        RECT  0.990 3.450 1.230 4.180 ;
        RECT  0.750 2.250 1.030 2.490 ;
        RECT  0.750 3.450 0.990 3.690 ;
        RECT  0.510 2.250 0.750 3.690 ;
    END
END ADDHX2

MACRO ADDHX1
    CLASS CORE ;
    FOREIGN ADDHX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ ADDHXL ;
    SIZE 8.580 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  3.500 2.950 3.510 3.220 ;
        RECT  3.510 2.950 3.750 3.520 ;
        RECT  3.570 1.190 3.810 1.620 ;
        RECT  3.750 2.950 4.470 3.220 ;
        RECT  3.810 1.380 4.470 1.620 ;
        RECT  4.470 1.380 4.710 3.220 ;
        RECT  4.710 2.950 4.720 3.220 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  7.460 1.270 7.810 1.530 ;
        RECT  7.810 1.260 8.010 1.540 ;
        RECT  8.010 1.230 8.130 1.630 ;
        RECT  8.010 2.970 8.170 3.370 ;
        RECT  8.130 1.230 8.170 1.840 ;
        RECT  8.170 1.230 8.410 3.370 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  1.840 2.430 2.240 2.830 ;
        RECT  2.240 2.430 2.750 2.750 ;
        RECT  2.750 2.430 2.990 3.220 ;
        RECT  2.990 2.430 3.230 4.250 ;
        RECT  3.230 2.430 3.600 2.670 ;
        RECT  3.600 1.900 3.840 2.670 ;
        RECT  3.840 1.900 4.190 2.140 ;
        RECT  3.230 4.010 5.510 4.250 ;
        RECT  5.510 3.350 5.750 4.250 ;
        RECT  5.750 3.350 6.650 3.590 ;
        RECT  6.650 3.180 6.890 3.590 ;
        RECT  6.890 3.180 7.050 3.580 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.950 1.830 5.850 2.230 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 4.480 1.390 5.440 ;
        RECT  1.390 4.640 6.970 5.440 ;
        RECT  6.970 4.480 7.950 5.440 ;
        RECT  7.950 4.640 8.580 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        RECT  0.990 -0.400 1.390 0.560 ;
        RECT  1.390 -0.400 5.070 0.400 ;
        RECT  5.070 -0.400 5.470 0.560 ;
        RECT  5.470 -0.400 7.900 0.400 ;
        RECT  7.900 -0.400 8.300 0.560 ;
        RECT  8.300 -0.400 8.580 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  7.730 1.950 7.880 2.350 ;
        RECT  7.490 1.950 7.730 4.110 ;
        RECT  7.480 1.950 7.490 2.350 ;
        RECT  6.100 3.870 7.490 4.110 ;
        RECT  7.080 1.960 7.480 2.200 ;
        RECT  6.840 0.640 7.080 2.200 ;
        RECT  6.650 0.640 6.840 0.880 ;
        RECT  6.130 1.310 6.370 3.070 ;
        RECT  5.360 1.310 6.130 1.550 ;
        RECT  5.230 2.830 6.130 3.070 ;
        RECT  5.120 0.860 5.360 1.550 ;
        RECT  4.990 2.830 5.230 3.730 ;
        RECT  4.650 0.860 5.120 1.100 ;
        RECT  4.190 3.490 4.990 3.730 ;
        RECT  4.250 0.670 4.650 1.100 ;
        RECT  3.290 0.670 4.250 0.910 ;
        RECT  3.050 0.670 3.290 2.140 ;
        RECT  1.440 1.900 3.050 2.140 ;
        RECT  2.530 0.700 2.770 1.100 ;
        RECT  2.470 3.640 2.710 4.180 ;
        RECT  0.920 1.380 2.680 1.620 ;
        RECT  0.570 0.860 2.530 1.100 ;
        RECT  0.570 3.940 2.470 4.180 ;
        RECT  1.540 3.380 2.050 3.620 ;
        RECT  1.300 2.980 1.540 3.620 ;
        RECT  1.200 1.900 1.440 2.700 ;
        RECT  0.920 2.980 1.300 3.220 ;
        RECT  0.680 1.380 0.920 3.220 ;
        RECT  0.400 0.700 0.570 1.100 ;
        RECT  0.400 3.500 0.570 4.180 ;
        RECT  0.160 0.700 0.400 4.180 ;
    END
END ADDHX1

MACRO ADDFHXL
    CLASS CORE ;
    FOREIGN ADDFHXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.720 1.830 14.830 2.090 ;
        RECT  14.830 1.820 15.270 2.090 ;
        RECT  15.270 3.050 15.430 3.450 ;
        RECT  15.270 1.390 15.430 2.090 ;
        RECT  15.430 1.390 15.670 3.450 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.620 2.960 13.730 3.360 ;
        RECT  13.730 1.380 13.970 3.360 ;
        RECT  13.970 2.950 14.020 3.360 ;
        RECT  13.970 1.380 14.130 1.780 ;
        RECT  14.020 2.950 14.320 3.210 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  12.650 2.370 13.100 2.790 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  6.800 2.950 6.970 3.210 ;
        RECT  6.970 2.640 7.060 3.210 ;
        RECT  7.060 2.640 7.290 3.200 ;
        RECT  7.290 2.640 7.370 3.040 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.860 2.390 0.900 2.650 ;
        RECT  0.900 2.140 1.120 2.650 ;
        RECT  1.120 2.140 1.300 2.640 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 1.330 5.440 ;
        RECT  1.330 3.980 1.340 5.440 ;
        RECT  1.340 3.780 1.740 5.440 ;
        RECT  1.740 3.980 1.750 5.440 ;
        RECT  1.750 4.640 6.820 5.440 ;
        RECT  6.820 4.480 7.220 5.440 ;
        RECT  7.220 4.640 11.380 5.440 ;
        RECT  11.380 4.480 12.360 5.440 ;
        RECT  12.360 4.640 14.450 5.440 ;
        RECT  14.450 4.480 14.850 5.440 ;
        RECT  14.850 4.640 15.840 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.090 0.400 ;
        RECT  1.090 -0.400 1.490 0.560 ;
        RECT  1.490 -0.400 7.820 0.400 ;
        RECT  7.820 -0.400 8.220 0.560 ;
        RECT  8.220 -0.400 12.220 0.400 ;
        RECT  12.220 -0.400 12.620 0.560 ;
        RECT  12.620 -0.400 14.610 0.400 ;
        RECT  14.610 -0.400 15.010 0.560 ;
        RECT  15.010 -0.400 15.840 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.990 2.370 15.150 2.770 ;
        RECT  14.750 2.370 14.990 4.180 ;
        RECT  10.540 3.940 14.750 4.180 ;
        RECT  9.640 0.860 14.370 1.100 ;
        RECT  12.990 1.380 13.390 1.780 ;
        RECT  12.830 3.170 13.230 3.570 ;
        RECT  12.380 1.380 12.990 1.620 ;
        RECT  12.380 3.170 12.830 3.410 ;
        RECT  12.140 1.380 12.380 3.410 ;
        RECT  10.210 1.380 12.140 1.620 ;
        RECT  11.890 2.610 12.140 3.010 ;
        RECT  11.610 1.900 11.810 2.140 ;
        RECT  11.370 1.900 11.610 3.500 ;
        RECT  11.220 3.260 11.370 3.500 ;
        RECT  10.820 3.260 11.220 3.660 ;
        RECT  10.970 1.900 11.050 2.140 ;
        RECT  10.730 1.900 10.970 2.980 ;
        RECT  10.650 1.900 10.730 2.140 ;
        RECT  10.540 2.740 10.730 2.980 ;
        RECT  10.300 2.740 10.540 4.180 ;
        RECT  10.060 3.340 10.300 3.740 ;
        RECT  9.970 1.380 10.210 2.460 ;
        RECT  9.780 2.220 9.970 2.460 ;
        RECT  9.540 2.220 9.780 3.690 ;
        RECT  9.420 0.860 9.640 1.780 ;
        RECT  9.380 3.290 9.540 3.690 ;
        RECT  9.400 0.860 9.420 1.940 ;
        RECT  9.260 1.540 9.400 1.940 ;
        RECT  9.100 1.540 9.260 2.980 ;
        RECT  8.740 0.680 9.120 1.100 ;
        RECT  9.020 1.540 9.100 3.890 ;
        RECT  8.860 2.740 9.020 3.890 ;
        RECT  8.460 3.650 8.860 3.890 ;
        RECT  8.720 0.680 8.740 2.460 ;
        RECT  8.580 0.860 8.720 2.460 ;
        RECT  8.500 0.860 8.580 3.040 ;
        RECT  7.420 0.860 8.500 1.100 ;
        RECT  8.340 2.220 8.500 3.040 ;
        RECT  8.060 1.540 8.220 1.940 ;
        RECT  8.060 3.390 8.100 3.790 ;
        RECT  7.820 1.540 8.060 3.790 ;
        RECT  7.700 3.390 7.820 3.790 ;
        RECT  6.380 3.490 7.700 3.730 ;
        RECT  7.300 1.890 7.540 2.290 ;
        RECT  7.180 0.670 7.420 1.100 ;
        RECT  6.900 1.890 7.300 2.130 ;
        RECT  4.820 0.670 7.180 0.910 ;
        RECT  6.660 1.190 6.900 2.130 ;
        RECT  5.340 1.190 6.660 1.430 ;
        RECT  6.140 2.230 6.380 3.730 ;
        RECT  5.860 1.710 6.260 1.950 ;
        RECT  5.620 1.710 5.860 4.210 ;
        RECT  2.670 3.970 5.620 4.210 ;
        RECT  5.100 1.190 5.340 3.690 ;
        RECT  3.440 3.450 5.100 3.690 ;
        RECT  4.580 0.670 4.820 3.170 ;
        RECT  4.060 1.090 4.140 1.490 ;
        RECT  4.060 2.770 4.140 3.170 ;
        RECT  3.980 1.090 4.060 3.170 ;
        RECT  3.820 0.680 3.980 3.170 ;
        RECT  3.740 0.680 3.820 1.490 ;
        RECT  3.740 2.770 3.820 3.170 ;
        RECT  2.010 0.680 3.740 0.920 ;
        RECT  3.200 1.270 3.440 3.690 ;
        RECT  2.980 1.270 3.200 1.510 ;
        RECT  2.980 3.150 3.200 3.690 ;
        RECT  2.430 1.200 2.670 4.210 ;
        RECT  2.290 1.200 2.430 1.600 ;
        RECT  2.220 3.240 2.430 3.640 ;
        RECT  1.880 2.200 2.040 2.600 ;
        RECT  1.770 0.680 2.010 1.100 ;
        RECT  1.640 1.550 1.880 3.170 ;
        RECT  0.610 0.860 1.770 1.100 ;
        RECT  0.920 1.550 1.640 1.790 ;
        RECT  0.920 2.930 1.640 3.170 ;
        RECT  0.680 1.390 0.920 1.790 ;
        RECT  0.680 2.930 0.920 3.330 ;
        RECT  0.460 3.740 0.860 4.140 ;
        RECT  0.400 0.670 0.610 1.100 ;
        RECT  0.400 3.740 0.460 3.980 ;
        RECT  0.160 0.670 0.400 3.980 ;
    END
END ADDFHXL

MACRO ADDFHX4
    CLASS CORE ;
    FOREIGN ADDFHX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ ADDFHXL ;
    SIZE 24.420 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  23.210 1.820 23.220 3.220 ;
        RECT  23.220 1.320 23.240 3.220 ;
        RECT  23.240 1.320 23.620 3.290 ;
        RECT  23.620 1.820 23.640 3.290 ;
        RECT  23.640 1.820 23.650 3.220 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.700 2.890 21.890 3.290 ;
        RECT  21.880 1.320 21.890 2.220 ;
        RECT  21.890 1.320 21.900 3.290 ;
        RECT  21.900 1.320 22.280 3.300 ;
        RECT  22.280 1.820 22.330 3.300 ;
        RECT  22.330 2.310 22.340 3.300 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  20.020 2.180 20.660 2.580 ;
        RECT  20.660 2.180 20.920 2.650 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  13.750 2.680 14.720 3.080 ;
        RECT  14.720 2.680 14.980 3.210 ;
        RECT  14.980 2.680 15.290 3.080 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.770 2.180 1.240 2.660 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.920 5.440 ;
        RECT  0.920 4.210 0.930 5.440 ;
        RECT  0.930 4.010 1.330 5.440 ;
        RECT  1.330 4.210 1.340 5.440 ;
        RECT  1.340 4.640 3.200 5.440 ;
        RECT  3.200 3.730 3.210 5.440 ;
        RECT  3.210 3.530 3.610 5.440 ;
        RECT  3.610 3.730 3.620 5.440 ;
        RECT  3.620 4.640 13.280 5.440 ;
        RECT  13.280 4.210 13.290 5.440 ;
        RECT  13.290 4.010 13.690 5.440 ;
        RECT  13.690 4.210 13.700 5.440 ;
        RECT  13.700 4.640 14.800 5.440 ;
        RECT  14.800 4.210 14.810 5.440 ;
        RECT  14.810 4.010 15.210 5.440 ;
        RECT  15.210 4.210 15.220 5.440 ;
        RECT  15.220 4.640 19.310 5.440 ;
        RECT  19.310 4.480 19.710 5.440 ;
        RECT  19.710 4.640 21.000 5.440 ;
        RECT  21.000 4.480 21.400 5.440 ;
        RECT  21.400 4.640 22.460 5.440 ;
        RECT  22.460 4.350 22.470 5.440 ;
        RECT  22.470 4.150 22.870 5.440 ;
        RECT  22.870 4.350 22.880 5.440 ;
        RECT  22.880 4.640 23.850 5.440 ;
        RECT  23.850 4.370 23.860 5.440 ;
        RECT  23.860 4.170 24.260 5.440 ;
        RECT  24.260 4.370 24.270 5.440 ;
        RECT  24.270 4.640 24.420 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        RECT  0.780 -0.400 1.180 0.560 ;
        RECT  1.180 -0.400 3.020 0.400 ;
        RECT  3.020 -0.400 3.420 0.560 ;
        RECT  3.420 -0.400 14.090 0.400 ;
        RECT  14.090 -0.400 14.490 0.560 ;
        RECT  14.490 -0.400 20.520 0.400 ;
        RECT  20.520 -0.400 21.500 0.560 ;
        RECT  21.500 -0.400 22.540 0.400 ;
        RECT  22.540 -0.400 22.550 0.840 ;
        RECT  22.550 -0.400 22.950 1.040 ;
        RECT  22.950 -0.400 22.960 0.840 ;
        RECT  22.960 -0.400 23.860 0.400 ;
        RECT  23.860 -0.400 24.260 1.040 ;
        RECT  24.260 -0.400 24.420 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  23.890 2.180 24.130 3.810 ;
        RECT  21.250 3.570 23.890 3.810 ;
        RECT  21.400 0.860 21.640 2.650 ;
        RECT  20.280 0.860 21.400 1.100 ;
        RECT  21.010 3.570 21.250 4.180 ;
        RECT  18.190 3.940 21.010 4.180 ;
        RECT  19.750 1.380 20.750 1.620 ;
        RECT  20.200 3.260 20.600 3.660 ;
        RECT  20.040 0.680 20.280 1.100 ;
        RECT  19.530 3.260 20.200 3.500 ;
        RECT  16.840 0.680 20.040 0.920 ;
        RECT  19.530 1.200 19.750 2.540 ;
        RECT  19.510 1.200 19.530 3.500 ;
        RECT  17.390 1.200 19.510 1.440 ;
        RECT  19.290 2.300 19.510 3.500 ;
        RECT  19.050 1.720 19.270 1.960 ;
        RECT  18.810 1.720 19.050 3.400 ;
        RECT  18.510 3.000 18.810 3.400 ;
        RECT  18.120 1.720 18.530 1.960 ;
        RECT  18.120 3.210 18.190 4.190 ;
        RECT  17.880 1.720 18.120 4.190 ;
        RECT  17.790 3.210 17.880 4.190 ;
        RECT  17.150 1.200 17.390 4.050 ;
        RECT  16.600 0.680 16.840 3.730 ;
        RECT  16.330 3.330 16.600 3.730 ;
        RECT  16.080 0.670 16.320 2.900 ;
        RECT  15.850 0.670 16.080 1.100 ;
        RECT  15.800 3.400 15.970 3.800 ;
        RECT  12.550 0.860 15.850 1.100 ;
        RECT  15.570 1.380 15.800 3.800 ;
        RECT  15.560 1.380 15.570 3.730 ;
        RECT  14.760 1.380 15.560 1.620 ;
        RECT  14.450 3.490 15.560 3.730 ;
        RECT  15.040 1.900 15.280 2.300 ;
        RECT  14.260 1.900 15.040 2.140 ;
        RECT  14.050 3.490 14.450 3.890 ;
        RECT  14.020 1.380 14.260 2.140 ;
        RECT  13.160 3.490 14.050 3.730 ;
        RECT  12.030 1.380 14.020 1.620 ;
        RECT  13.160 1.900 13.730 2.140 ;
        RECT  12.920 1.900 13.160 3.730 ;
        RECT  12.840 1.900 12.920 3.520 ;
        RECT  12.320 1.930 12.560 4.360 ;
        RECT  12.310 0.680 12.550 1.100 ;
        RECT  11.510 1.930 12.320 2.170 ;
        RECT  10.620 4.120 12.320 4.360 ;
        RECT  10.310 0.680 12.310 0.920 ;
        RECT  11.800 2.450 12.040 3.840 ;
        RECT  11.790 1.200 12.030 1.620 ;
        RECT  10.830 2.450 11.800 2.690 ;
        RECT  10.020 3.600 11.800 3.840 ;
        RECT  10.830 1.200 11.790 1.440 ;
        RECT  10.310 3.080 11.520 3.320 ;
        RECT  11.110 1.720 11.510 2.170 ;
        RECT  10.590 1.200 10.830 2.690 ;
        RECT  10.300 4.120 10.620 4.370 ;
        RECT  10.070 0.670 10.310 3.320 ;
        RECT  4.370 4.130 10.300 4.370 ;
        RECT  8.740 0.670 10.070 0.910 ;
        RECT  9.780 3.600 10.020 3.850 ;
        RECT  7.390 3.610 9.780 3.850 ;
        RECT  9.500 2.860 9.710 3.260 ;
        RECT  9.260 1.190 9.500 3.330 ;
        RECT  9.100 1.190 9.260 1.430 ;
        RECT  7.990 3.090 9.260 3.330 ;
        RECT  8.740 2.570 8.970 2.810 ;
        RECT  8.500 0.670 8.740 2.810 ;
        RECT  8.340 0.960 8.500 1.360 ;
        RECT  7.980 1.040 7.990 3.330 ;
        RECT  7.820 0.960 7.980 3.330 ;
        RECT  7.750 0.670 7.820 3.330 ;
        RECT  7.580 0.670 7.750 1.360 ;
        RECT  6.480 0.670 7.580 0.910 ;
        RECT  7.230 3.280 7.390 3.850 ;
        RECT  6.990 1.190 7.230 3.850 ;
        RECT  6.820 1.190 6.990 1.430 ;
        RECT  5.130 3.610 6.990 3.850 ;
        RECT  6.480 3.080 6.630 3.320 ;
        RECT  6.240 0.670 6.480 3.320 ;
        RECT  6.000 0.670 6.240 1.070 ;
        RECT  6.230 3.080 6.240 3.320 ;
        RECT  3.940 0.680 6.000 0.920 ;
        RECT  5.660 1.410 5.900 1.810 ;
        RECT  5.660 3.080 5.890 3.320 ;
        RECT  5.420 1.200 5.660 3.320 ;
        RECT  4.460 1.200 5.420 1.440 ;
        RECT  4.980 1.720 5.140 1.960 ;
        RECT  4.980 3.000 5.130 3.850 ;
        RECT  4.890 1.720 4.980 3.850 ;
        RECT  4.740 1.720 4.890 3.400 ;
        RECT  4.730 3.000 4.740 3.400 ;
        RECT  4.340 1.200 4.460 1.780 ;
        RECT  4.340 3.000 4.370 4.370 ;
        RECT  4.220 1.200 4.340 4.370 ;
        RECT  4.130 1.380 4.220 4.370 ;
        RECT  4.100 1.380 4.130 3.530 ;
        RECT  3.980 1.380 4.100 1.780 ;
        RECT  3.970 3.000 4.100 3.530 ;
        RECT  2.740 1.380 3.980 1.620 ;
        RECT  2.870 3.000 3.970 3.240 ;
        RECT  3.700 0.680 3.940 1.100 ;
        RECT  2.850 2.060 3.830 2.460 ;
        RECT  0.660 0.860 3.700 1.100 ;
        RECT  2.470 3.000 2.870 4.020 ;
        RECT  2.130 2.060 2.850 2.300 ;
        RECT  2.340 1.380 2.740 1.780 ;
        RECT  2.000 2.060 2.130 3.210 ;
        RECT  1.950 4.070 2.110 4.310 ;
        RECT  1.760 1.380 2.000 3.210 ;
        RECT  1.710 3.490 1.950 4.310 ;
        RECT  1.600 1.380 1.760 1.780 ;
        RECT  1.750 2.220 1.760 3.210 ;
        RECT  1.730 2.810 1.750 3.210 ;
        RECT  0.570 3.490 1.710 3.730 ;
        RECT  0.500 0.860 0.660 1.790 ;
        RECT  0.500 2.960 0.570 3.940 ;
        RECT  0.420 0.860 0.500 3.940 ;
        RECT  0.260 1.390 0.420 3.940 ;
        RECT  0.170 2.960 0.260 3.940 ;
    END
END ADDFHX4

MACRO ADDFHX2
    CLASS CORE ;
    FOREIGN ADDFHX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ ADDFHXL ;
    SIZE 24.420 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  23.840 1.550 23.850 1.860 ;
        RECT  23.850 0.720 23.960 1.860 ;
        RECT  23.850 3.030 23.980 4.010 ;
        RECT  23.960 0.720 23.980 2.090 ;
        RECT  23.980 0.720 24.220 4.010 ;
        RECT  24.220 3.030 24.250 4.010 ;
        RECT  24.220 0.720 24.250 1.860 ;
        RECT  24.250 1.390 24.260 1.860 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  21.980 2.950 22.310 3.210 ;
        RECT  22.310 2.830 22.470 3.230 ;
        RECT  22.370 1.380 22.470 1.780 ;
        RECT  22.470 1.380 22.710 3.230 ;
        RECT  22.710 1.380 22.770 1.840 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  20.470 2.320 21.450 2.720 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  14.050 2.640 14.720 3.040 ;
        RECT  14.720 2.640 14.980 3.210 ;
        RECT  14.980 2.640 15.590 3.040 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.820 2.180 1.240 2.660 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.920 5.440 ;
        RECT  0.920 4.210 0.930 5.440 ;
        RECT  0.930 4.010 1.330 5.440 ;
        RECT  1.330 4.210 1.340 5.440 ;
        RECT  1.340 4.640 3.200 5.440 ;
        RECT  3.200 3.730 3.210 5.440 ;
        RECT  3.210 3.530 3.610 5.440 ;
        RECT  3.610 3.730 3.620 5.440 ;
        RECT  3.620 4.640 13.580 5.440 ;
        RECT  13.580 4.210 13.590 5.440 ;
        RECT  13.590 4.010 13.990 5.440 ;
        RECT  13.990 4.210 14.000 5.440 ;
        RECT  14.000 4.640 15.100 5.440 ;
        RECT  15.100 4.210 15.110 5.440 ;
        RECT  15.110 4.010 15.510 5.440 ;
        RECT  15.510 4.210 15.520 5.440 ;
        RECT  15.520 4.640 19.730 5.440 ;
        RECT  19.730 4.480 20.130 5.440 ;
        RECT  20.130 4.640 21.490 5.440 ;
        RECT  21.490 4.480 21.890 5.440 ;
        RECT  21.890 4.640 23.010 5.440 ;
        RECT  23.010 4.030 23.410 5.440 ;
        RECT  23.410 4.640 24.420 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.780 0.400 ;
        RECT  0.780 -0.400 1.180 0.560 ;
        RECT  1.180 -0.400 3.020 0.400 ;
        RECT  3.020 -0.400 3.420 0.560 ;
        RECT  3.420 -0.400 14.210 0.400 ;
        RECT  14.210 -0.400 14.610 0.560 ;
        RECT  14.610 -0.400 20.980 0.400 ;
        RECT  20.980 -0.400 21.960 0.560 ;
        RECT  21.960 -0.400 23.090 0.400 ;
        RECT  23.090 -0.400 23.490 1.040 ;
        RECT  23.490 -0.400 24.420 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  23.430 2.260 23.590 2.660 ;
        RECT  23.190 2.260 23.430 3.750 ;
        RECT  21.590 3.510 23.190 3.750 ;
        RECT  22.030 2.060 22.190 2.460 ;
        RECT  21.790 0.860 22.030 2.460 ;
        RECT  20.710 0.860 21.790 1.100 ;
        RECT  21.350 3.510 21.590 4.180 ;
        RECT  18.550 3.940 21.350 4.180 ;
        RECT  20.800 1.380 21.200 1.780 ;
        RECT  20.670 3.260 21.070 3.660 ;
        RECT  20.190 1.460 20.800 1.700 ;
        RECT  20.470 0.680 20.710 1.100 ;
        RECT  20.190 3.260 20.670 3.500 ;
        RECT  17.140 0.680 20.470 0.920 ;
        RECT  19.950 1.200 20.190 3.500 ;
        RECT  17.710 1.200 19.950 1.440 ;
        RECT  19.710 2.300 19.950 2.700 ;
        RECT  19.430 1.720 19.670 1.960 ;
        RECT  19.190 1.720 19.430 3.400 ;
        RECT  18.910 3.000 19.190 3.400 ;
        RECT  18.460 1.720 18.910 1.960 ;
        RECT  18.460 3.210 18.550 4.190 ;
        RECT  18.220 1.720 18.460 4.190 ;
        RECT  18.150 3.210 18.220 4.190 ;
        RECT  17.470 1.200 17.710 4.050 ;
        RECT  16.900 0.680 17.140 3.730 ;
        RECT  16.630 3.330 16.900 3.730 ;
        RECT  16.380 0.670 16.620 2.900 ;
        RECT  16.120 0.670 16.380 1.100 ;
        RECT  16.100 3.400 16.270 3.800 ;
        RECT  12.550 0.860 16.120 1.100 ;
        RECT  15.870 1.380 16.100 3.800 ;
        RECT  15.860 1.380 15.870 3.730 ;
        RECT  15.030 1.380 15.860 1.620 ;
        RECT  14.750 3.490 15.860 3.730 ;
        RECT  15.310 1.900 15.550 2.320 ;
        RECT  14.620 1.900 15.310 2.140 ;
        RECT  14.350 3.490 14.750 3.890 ;
        RECT  14.380 1.380 14.620 2.140 ;
        RECT  12.030 1.380 14.380 1.620 ;
        RECT  13.080 3.490 14.350 3.730 ;
        RECT  13.080 1.900 13.730 2.140 ;
        RECT  12.840 1.900 13.080 3.730 ;
        RECT  12.320 1.930 12.560 4.350 ;
        RECT  12.310 0.670 12.550 1.100 ;
        RECT  11.510 1.930 12.320 2.170 ;
        RECT  10.620 4.110 12.320 4.350 ;
        RECT  10.310 0.670 12.310 0.910 ;
        RECT  11.800 2.450 12.040 3.830 ;
        RECT  11.790 1.190 12.030 1.620 ;
        RECT  10.830 2.450 11.800 2.690 ;
        RECT  10.020 3.590 11.800 3.830 ;
        RECT  10.830 1.190 11.790 1.430 ;
        RECT  10.310 3.070 11.520 3.310 ;
        RECT  11.110 1.710 11.510 2.170 ;
        RECT  10.590 1.190 10.830 2.690 ;
        RECT  10.300 4.110 10.620 4.370 ;
        RECT  10.070 0.670 10.310 3.310 ;
        RECT  4.370 4.130 10.300 4.370 ;
        RECT  8.740 0.670 10.070 0.910 ;
        RECT  9.780 3.590 10.020 3.850 ;
        RECT  7.390 3.610 9.780 3.850 ;
        RECT  9.500 2.860 9.710 3.260 ;
        RECT  9.260 1.190 9.500 3.330 ;
        RECT  9.100 1.190 9.260 1.430 ;
        RECT  7.990 3.090 9.260 3.330 ;
        RECT  8.740 2.570 8.970 2.810 ;
        RECT  8.500 0.670 8.740 2.810 ;
        RECT  8.340 0.960 8.500 1.360 ;
        RECT  7.980 1.040 7.990 3.330 ;
        RECT  7.820 0.960 7.980 3.330 ;
        RECT  7.750 0.670 7.820 3.330 ;
        RECT  7.580 0.670 7.750 1.360 ;
        RECT  6.480 0.670 7.580 0.910 ;
        RECT  7.230 3.280 7.390 3.850 ;
        RECT  6.990 1.190 7.230 3.850 ;
        RECT  6.820 1.190 6.990 1.430 ;
        RECT  5.130 3.610 6.990 3.850 ;
        RECT  6.480 3.080 6.630 3.320 ;
        RECT  6.240 0.670 6.480 3.320 ;
        RECT  6.000 0.670 6.240 1.070 ;
        RECT  6.230 3.080 6.240 3.320 ;
        RECT  3.940 0.680 6.000 0.920 ;
        RECT  5.660 1.410 5.900 1.810 ;
        RECT  5.660 3.080 5.890 3.320 ;
        RECT  5.420 1.200 5.660 3.320 ;
        RECT  4.460 1.200 5.420 1.440 ;
        RECT  4.980 1.720 5.140 1.960 ;
        RECT  4.980 3.000 5.130 3.850 ;
        RECT  4.890 1.720 4.980 3.850 ;
        RECT  4.740 1.720 4.890 3.400 ;
        RECT  4.730 3.000 4.740 3.400 ;
        RECT  4.340 1.200 4.460 1.780 ;
        RECT  4.340 3.000 4.370 4.370 ;
        RECT  4.220 1.200 4.340 4.370 ;
        RECT  4.130 1.380 4.220 4.370 ;
        RECT  4.100 1.380 4.130 3.530 ;
        RECT  3.980 1.380 4.100 1.780 ;
        RECT  3.970 3.000 4.100 3.530 ;
        RECT  2.740 1.380 3.980 1.620 ;
        RECT  2.850 3.000 3.970 3.240 ;
        RECT  3.700 0.680 3.940 1.100 ;
        RECT  2.850 2.060 3.830 2.460 ;
        RECT  0.660 0.860 3.700 1.100 ;
        RECT  2.110 2.060 2.850 2.300 ;
        RECT  2.450 2.990 2.850 3.950 ;
        RECT  2.340 1.380 2.740 1.780 ;
        RECT  2.000 2.060 2.110 3.210 ;
        RECT  1.950 4.070 2.110 4.310 ;
        RECT  1.870 1.380 2.000 3.210 ;
        RECT  1.710 3.490 1.950 4.310 ;
        RECT  1.760 1.380 1.870 2.300 ;
        RECT  1.710 2.810 1.870 3.210 ;
        RECT  1.720 1.380 1.760 2.110 ;
        RECT  1.600 1.380 1.720 1.780 ;
        RECT  0.570 3.490 1.710 3.730 ;
        RECT  0.500 0.860 0.660 1.790 ;
        RECT  0.500 2.960 0.570 3.940 ;
        RECT  0.420 0.860 0.500 3.940 ;
        RECT  0.260 1.390 0.420 3.940 ;
        RECT  0.170 2.960 0.260 3.940 ;
    END
END ADDFHX2

MACRO ADDFHX1
    CLASS CORE ;
    FOREIGN ADDFHX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ ADDFHXL ;
    SIZE 17.160 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  16.040 1.270 16.300 1.540 ;
        RECT  16.300 1.300 16.590 1.540 ;
        RECT  16.590 1.300 16.610 1.720 ;
        RECT  16.590 3.130 16.660 3.530 ;
        RECT  16.610 1.300 16.660 1.820 ;
        RECT  16.660 1.300 16.900 3.530 ;
        RECT  16.900 3.130 16.990 3.530 ;
        RECT  16.900 1.320 16.990 1.840 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.720 2.950 14.730 3.210 ;
        RECT  14.730 2.950 14.950 3.540 ;
        RECT  14.950 1.380 15.190 3.540 ;
        RECT  15.190 3.140 15.250 3.540 ;
        RECT  15.190 1.380 15.350 1.780 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  13.790 2.380 13.990 2.780 ;
        RECT  13.990 2.370 14.320 2.790 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  7.620 2.210 8.020 3.190 ;
        RECT  8.020 2.940 8.030 3.190 ;
        RECT  8.030 2.950 8.120 3.190 ;
        RECT  8.120 2.950 8.380 3.210 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.790 1.990 0.860 2.390 ;
        RECT  0.860 1.830 1.120 2.390 ;
        RECT  1.120 1.990 1.190 2.390 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.930 5.440 ;
        RECT  0.930 2.750 1.330 5.440 ;
        RECT  1.330 4.640 2.220 5.440 ;
        RECT  2.220 3.700 2.230 5.440 ;
        RECT  2.230 3.500 2.630 5.440 ;
        RECT  2.630 3.700 2.640 5.440 ;
        RECT  2.640 4.640 7.730 5.440 ;
        RECT  7.730 4.480 8.130 5.440 ;
        RECT  8.130 4.640 12.500 5.440 ;
        RECT  12.500 4.480 13.480 5.440 ;
        RECT  13.480 4.640 15.680 5.440 ;
        RECT  15.680 4.480 16.080 5.440 ;
        RECT  16.080 4.640 17.160 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.020 0.400 ;
        RECT  1.020 -0.400 2.000 0.560 ;
        RECT  2.000 -0.400 8.350 0.400 ;
        RECT  8.350 -0.400 8.750 0.560 ;
        RECT  8.750 -0.400 13.390 0.400 ;
        RECT  13.390 -0.400 13.790 0.560 ;
        RECT  13.790 -0.400 15.770 0.400 ;
        RECT  15.770 -0.400 16.170 0.560 ;
        RECT  16.170 -0.400 17.160 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  16.260 2.350 16.420 2.750 ;
        RECT  16.020 2.350 16.260 4.180 ;
        RECT  11.580 3.940 16.020 4.180 ;
        RECT  15.090 0.680 15.490 1.100 ;
        RECT  10.460 0.860 15.090 1.100 ;
        RECT  14.200 1.380 14.600 1.780 ;
        RECT  13.890 3.190 14.290 3.590 ;
        RECT  13.510 1.380 14.200 1.620 ;
        RECT  13.510 3.190 13.890 3.430 ;
        RECT  13.270 1.380 13.510 3.430 ;
        RECT  11.360 1.380 13.270 1.620 ;
        RECT  13.010 2.610 13.270 3.010 ;
        RECT  12.730 1.900 12.970 2.140 ;
        RECT  12.490 1.900 12.730 3.420 ;
        RECT  12.340 3.180 12.490 3.420 ;
        RECT  11.940 3.180 12.340 3.580 ;
        RECT  12.130 1.900 12.210 2.140 ;
        RECT  11.810 1.900 12.130 2.150 ;
        RECT  11.580 1.910 11.810 2.150 ;
        RECT  11.340 1.910 11.580 4.180 ;
        RECT  11.040 1.380 11.360 1.630 ;
        RECT  11.180 3.340 11.340 3.740 ;
        RECT  10.980 1.390 11.040 1.630 ;
        RECT  10.740 1.390 10.980 2.500 ;
        RECT  10.500 2.260 10.740 3.690 ;
        RECT  10.220 0.860 10.460 1.950 ;
        RECT  9.980 1.540 10.220 4.350 ;
        RECT  9.370 4.110 9.980 4.350 ;
        RECT  9.280 0.680 9.940 0.920 ;
        RECT  9.460 1.540 9.700 3.830 ;
        RECT  8.950 3.590 9.460 3.830 ;
        RECT  9.180 0.680 9.280 1.100 ;
        RECT  9.030 0.680 9.180 3.310 ;
        RECT  8.940 0.860 9.030 3.310 ;
        RECT  8.550 3.590 8.950 3.990 ;
        RECT  8.070 0.860 8.940 1.100 ;
        RECT  8.750 3.070 8.940 3.310 ;
        RECT  8.420 1.430 8.660 2.670 ;
        RECT  7.310 3.750 8.550 3.990 ;
        RECT  7.550 1.430 8.420 1.670 ;
        RECT  7.830 0.670 8.070 1.100 ;
        RECT  5.660 0.670 7.830 0.910 ;
        RECT  7.310 1.190 7.550 1.670 ;
        RECT  6.180 1.190 7.310 1.430 ;
        RECT  7.220 3.660 7.310 4.060 ;
        RECT  6.980 2.230 7.220 4.060 ;
        RECT  6.700 1.710 7.030 1.950 ;
        RECT  6.910 3.660 6.980 4.060 ;
        RECT  6.630 1.710 6.700 2.350 ;
        RECT  6.460 1.710 6.630 4.210 ;
        RECT  6.390 2.110 6.460 4.210 ;
        RECT  3.440 3.970 6.390 4.210 ;
        RECT  6.110 1.190 6.180 1.830 ;
        RECT  5.940 1.190 6.110 3.690 ;
        RECT  5.870 1.590 5.940 3.690 ;
        RECT  4.210 3.450 5.870 3.690 ;
        RECT  5.590 0.670 5.660 1.310 ;
        RECT  5.350 0.670 5.590 3.170 ;
        RECT  4.830 1.110 4.980 1.510 ;
        RECT  4.830 2.770 4.910 3.170 ;
        RECT  4.820 1.110 4.830 3.170 ;
        RECT  4.590 0.670 4.820 3.170 ;
        RECT  4.580 0.670 4.590 1.510 ;
        RECT  4.510 2.770 4.590 3.170 ;
        RECT  2.520 0.670 4.580 0.910 ;
        RECT  3.970 1.190 4.210 3.690 ;
        RECT  3.810 1.190 3.970 1.590 ;
        RECT  3.750 3.290 3.970 3.690 ;
        RECT  3.440 1.190 3.450 1.590 ;
        RECT  3.200 1.190 3.440 4.210 ;
        RECT  3.050 1.190 3.200 1.590 ;
        RECT  2.990 3.500 3.200 3.900 ;
        RECT  2.130 2.010 2.870 2.410 ;
        RECT  2.280 0.670 2.520 1.100 ;
        RECT  0.490 0.860 2.280 1.100 ;
        RECT  1.890 1.390 2.130 3.150 ;
        RECT  1.710 1.390 1.890 1.790 ;
        RECT  1.730 2.750 1.890 3.150 ;
        RECT  0.490 2.800 0.570 3.780 ;
        RECT  0.250 0.860 0.490 3.780 ;
        RECT  0.170 2.800 0.250 3.780 ;
    END
END ADDFHX1

MACRO ADDFXL
    CLASS CORE ;
    FOREIGN ADDFXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.090 2.750 13.250 3.150 ;
        RECT  12.940 1.380 13.250 1.780 ;
        RECT  13.250 1.380 13.490 3.150 ;
        RECT  13.490 2.390 13.660 2.650 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.610 2.840 14.630 3.240 ;
        RECT  14.630 2.510 14.720 3.240 ;
        RECT  14.720 2.390 14.730 3.240 ;
        RECT  14.610 1.390 14.730 1.960 ;
        RECT  14.730 1.390 14.970 3.240 ;
        RECT  14.970 2.390 14.980 3.240 ;
        RECT  14.980 2.510 15.010 3.240 ;
        RECT  14.970 1.390 15.010 1.960 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.970 1.960 10.010 2.200 ;
        RECT  10.100 2.950 10.130 3.210 ;
        RECT  10.010 1.960 10.130 2.400 ;
        RECT  10.130 1.960 10.370 3.440 ;
        RECT  10.370 2.960 10.630 3.440 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.210 2.090 ;
        RECT  0.210 1.830 0.460 2.420 ;
        RECT  0.460 2.010 0.700 2.420 ;
        RECT  0.700 2.010 0.810 2.410 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.630 2.320 5.170 2.720 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 4.480 1.390 5.440 ;
        RECT  1.390 4.640 9.920 5.440 ;
        RECT  9.920 3.920 9.930 5.440 ;
        RECT  9.930 3.720 10.330 5.440 ;
        RECT  10.330 3.920 10.340 5.440 ;
        RECT  10.340 4.640 13.840 5.440 ;
        RECT  13.840 3.130 13.850 5.440 ;
        RECT  13.850 2.930 14.250 5.440 ;
        RECT  14.250 3.130 14.260 5.440 ;
        RECT  14.260 4.640 15.180 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 1.050 0.400 ;
        RECT  1.050 -0.400 1.450 0.560 ;
        RECT  1.450 -0.400 4.880 0.400 ;
        RECT  4.880 -0.400 4.890 0.730 ;
        RECT  4.890 -0.400 5.290 0.850 ;
        RECT  5.290 -0.400 5.300 0.730 ;
        RECT  5.300 -0.400 10.570 0.400 ;
        RECT  10.570 -0.400 10.970 0.560 ;
        RECT  10.970 -0.400 13.820 0.400 ;
        RECT  13.820 -0.400 14.220 0.560 ;
        RECT  14.220 -0.400 15.180 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  13.170 3.850 13.570 4.250 ;
        RECT  11.990 3.880 13.170 4.120 ;
        RECT  12.590 3.190 12.750 3.590 ;
        RECT  12.430 1.340 12.590 3.590 ;
        RECT  12.350 0.870 12.430 3.590 ;
        RECT  12.190 0.870 12.350 1.740 ;
        RECT  10.330 0.870 12.190 1.110 ;
        RECT  11.830 3.200 11.990 4.120 ;
        RECT  11.750 1.390 11.830 4.120 ;
        RECT  11.590 1.390 11.750 3.600 ;
        RECT  11.430 1.390 11.590 1.790 ;
        RECT  10.910 1.390 11.150 3.500 ;
        RECT  10.650 1.390 10.910 1.790 ;
        RECT  9.850 1.440 10.650 1.680 ;
        RECT  10.090 0.680 10.330 1.110 ;
        RECT  6.490 0.680 10.090 0.920 ;
        RECT  9.610 1.200 9.850 1.680 ;
        RECT  9.460 2.320 9.650 2.720 ;
        RECT  7.130 1.200 9.610 1.440 ;
        RECT  9.450 2.310 9.460 3.410 ;
        RECT  9.370 2.310 9.450 3.610 ;
        RECT  9.130 1.720 9.370 3.610 ;
        RECT  9.050 2.310 9.130 3.610 ;
        RECT  9.040 2.310 9.050 3.410 ;
        RECT  8.370 1.720 8.610 4.370 ;
        RECT  8.090 3.970 8.370 4.370 ;
        RECT  7.850 1.880 8.090 3.500 ;
        RECT  7.730 1.880 7.850 2.120 ;
        RECT  7.480 3.260 7.850 3.500 ;
        RECT  7.490 1.720 7.730 2.120 ;
        RECT  7.500 2.500 7.570 2.970 ;
        RECT  7.130 2.490 7.500 2.970 ;
        RECT  7.320 3.260 7.480 3.660 ;
        RECT  7.080 3.260 7.320 4.360 ;
        RECT  6.890 1.200 7.130 2.970 ;
        RECT  5.820 4.060 7.080 4.360 ;
        RECT  6.690 2.730 6.890 2.970 ;
        RECT  6.450 2.730 6.690 3.780 ;
        RECT  6.250 0.680 6.490 1.640 ;
        RECT  5.810 1.930 6.490 2.340 ;
        RECT  6.290 3.240 6.450 3.780 ;
        RECT  3.770 3.540 6.290 3.780 ;
        RECT  6.090 1.130 6.250 1.640 ;
        RECT  4.610 1.130 6.090 1.370 ;
        RECT  5.810 3.020 5.930 3.260 ;
        RECT  1.910 4.120 5.820 4.360 ;
        RECT  5.570 1.650 5.810 3.260 ;
        RECT  4.030 1.650 5.570 1.890 ;
        RECT  4.050 3.020 5.570 3.260 ;
        RECT  4.370 0.870 4.610 1.370 ;
        RECT  2.690 0.870 4.370 1.110 ;
        RECT  3.790 1.390 4.030 1.890 ;
        RECT  3.530 2.330 3.770 3.780 ;
        RECT  3.470 2.330 3.530 2.570 ;
        RECT  3.230 1.550 3.470 2.570 ;
        RECT  3.010 3.440 3.250 3.840 ;
        RECT  3.210 1.550 3.230 1.790 ;
        RECT  2.970 1.390 3.210 1.790 ;
        RECT  2.950 2.870 3.190 3.110 ;
        RECT  2.430 3.440 3.010 3.680 ;
        RECT  2.710 2.070 2.950 3.110 ;
        RECT  2.690 2.070 2.710 2.310 ;
        RECT  2.450 0.870 2.690 2.310 ;
        RECT  2.190 2.910 2.430 3.680 ;
        RECT  2.170 2.910 2.190 3.310 ;
        RECT  1.930 1.390 2.170 3.310 ;
        RECT  1.840 2.910 1.930 3.310 ;
        RECT  1.670 3.650 1.910 4.360 ;
        RECT  1.470 3.650 1.670 3.890 ;
        RECT  1.470 2.010 1.650 2.410 ;
        RECT  1.230 1.310 1.470 3.890 ;
        RECT  0.570 1.310 1.230 1.550 ;
        RECT  0.170 3.490 1.230 3.890 ;
        RECT  0.170 1.150 0.570 1.550 ;
    END
END ADDFXL

MACRO ADDFX4
    CLASS CORE ;
    FOREIGN ADDFX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ ADDFXL ;
    SIZE 15.840 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.630 1.820 14.640 3.220 ;
        RECT  14.640 1.380 14.650 3.220 ;
        RECT  14.650 1.380 15.040 3.230 ;
        RECT  15.040 1.820 15.050 3.230 ;
        RECT  15.050 1.820 15.070 3.220 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.650 1.820 12.690 3.220 ;
        RECT  12.690 1.380 13.090 3.230 ;
        RECT  13.090 2.830 13.510 3.230 ;
        RECT  13.090 1.380 13.700 1.780 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.840 1.960 10.050 4.190 ;
        RECT  10.050 1.960 10.080 4.350 ;
        RECT  10.080 1.960 10.370 2.200 ;
        RECT  10.080 3.950 10.450 4.350 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.220 2.090 ;
        RECT  0.220 1.830 0.460 2.420 ;
        RECT  0.460 2.010 0.700 2.420 ;
        RECT  0.700 2.010 0.810 2.410 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.280 2.320 5.260 2.720 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 4.480 1.390 5.440 ;
        RECT  1.390 4.640 9.180 5.440 ;
        RECT  9.180 4.070 9.600 5.440 ;
        RECT  9.600 4.640 12.480 5.440 ;
        RECT  12.480 4.310 12.490 5.440 ;
        RECT  12.490 4.110 12.890 5.440 ;
        RECT  12.890 4.310 12.900 5.440 ;
        RECT  12.900 4.640 13.870 5.440 ;
        RECT  13.870 4.290 13.880 5.440 ;
        RECT  13.880 4.090 14.280 5.440 ;
        RECT  14.280 4.290 14.290 5.440 ;
        RECT  14.290 4.640 15.260 5.440 ;
        RECT  15.260 4.290 15.270 5.440 ;
        RECT  15.270 4.090 15.670 5.440 ;
        RECT  15.670 4.290 15.680 5.440 ;
        RECT  15.680 4.640 15.840 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        RECT  0.990 -0.400 1.390 0.560 ;
        RECT  1.390 -0.400 4.880 0.400 ;
        RECT  4.880 -0.400 4.890 0.730 ;
        RECT  4.890 -0.400 5.290 0.850 ;
        RECT  5.290 -0.400 5.300 0.730 ;
        RECT  5.300 -0.400 10.700 0.400 ;
        RECT  10.700 -0.400 11.100 0.560 ;
        RECT  11.100 -0.400 12.650 0.400 ;
        RECT  12.650 -0.400 12.660 0.900 ;
        RECT  12.660 -0.400 13.060 1.100 ;
        RECT  13.060 -0.400 13.070 0.900 ;
        RECT  13.070 -0.400 13.960 0.400 ;
        RECT  13.960 -0.400 13.970 0.900 ;
        RECT  13.970 -0.400 14.370 1.100 ;
        RECT  14.370 -0.400 14.380 0.900 ;
        RECT  14.380 -0.400 15.270 0.400 ;
        RECT  15.270 -0.400 15.280 0.900 ;
        RECT  15.280 -0.400 15.680 1.100 ;
        RECT  15.680 -0.400 15.690 0.900 ;
        RECT  15.690 -0.400 15.840 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  15.310 2.120 15.550 3.810 ;
        RECT  13.330 3.570 15.310 3.810 ;
        RECT  13.880 2.830 14.280 3.330 ;
        RECT  13.090 3.570 13.330 3.830 ;
        RECT  11.510 3.590 13.090 3.830 ;
        RECT  12.230 0.870 12.390 3.310 ;
        RECT  12.150 0.680 12.230 3.310 ;
        RECT  11.830 0.680 12.150 1.110 ;
        RECT  11.750 3.070 12.150 3.310 ;
        RECT  11.750 1.460 11.910 1.860 ;
        RECT  10.400 0.870 11.830 1.110 ;
        RECT  11.510 1.460 11.750 2.310 ;
        RECT  11.270 2.070 11.510 3.830 ;
        RECT  10.960 3.180 11.270 3.580 ;
        RECT  10.850 1.390 11.040 1.830 ;
        RECT  10.610 1.390 10.850 2.940 ;
        RECT  9.880 1.390 10.610 1.630 ;
        RECT  10.560 2.700 10.610 2.940 ;
        RECT  10.320 2.700 10.560 3.600 ;
        RECT  10.160 0.680 10.400 1.110 ;
        RECT  6.610 0.680 10.160 0.920 ;
        RECT  9.640 1.200 9.880 1.630 ;
        RECT  7.200 1.200 9.640 1.440 ;
        RECT  9.370 2.330 9.600 2.730 ;
        RECT  9.290 1.720 9.370 2.730 ;
        RECT  9.130 1.720 9.290 3.600 ;
        RECT  8.890 2.330 9.130 3.600 ;
        RECT  8.530 1.720 8.610 2.120 ;
        RECT  8.470 1.720 8.530 3.450 ;
        RECT  8.370 1.720 8.470 4.360 ;
        RECT  8.290 1.800 8.370 4.360 ;
        RECT  8.230 3.130 8.290 4.360 ;
        RECT  7.960 3.960 8.230 4.360 ;
        RECT  7.750 1.880 7.990 3.410 ;
        RECT  7.730 1.880 7.750 2.120 ;
        RECT  7.450 3.170 7.750 3.410 ;
        RECT  7.490 1.720 7.730 2.120 ;
        RECT  7.200 2.480 7.510 2.890 ;
        RECT  7.290 3.170 7.450 3.570 ;
        RECT  7.050 3.170 7.290 4.360 ;
        RECT  6.960 1.200 7.200 2.890 ;
        RECT  5.820 4.050 7.050 4.360 ;
        RECT  6.680 2.650 6.960 2.890 ;
        RECT  5.870 1.930 6.680 2.330 ;
        RECT  6.520 2.650 6.680 3.510 ;
        RECT  6.370 0.680 6.610 1.590 ;
        RECT  6.440 2.650 6.520 3.770 ;
        RECT  6.280 3.110 6.440 3.770 ;
        RECT  6.210 1.130 6.370 1.590 ;
        RECT  3.770 3.530 6.280 3.770 ;
        RECT  4.610 1.130 6.210 1.370 ;
        RECT  5.870 3.010 5.930 3.250 ;
        RECT  5.630 1.650 5.870 3.250 ;
        RECT  1.910 4.120 5.820 4.360 ;
        RECT  4.090 1.650 5.630 1.890 ;
        RECT  4.050 3.010 5.630 3.250 ;
        RECT  4.370 0.870 4.610 1.370 ;
        RECT  2.690 0.870 4.370 1.110 ;
        RECT  3.850 1.390 4.090 1.890 ;
        RECT  3.530 2.330 3.770 3.770 ;
        RECT  3.470 2.330 3.530 2.570 ;
        RECT  3.230 1.550 3.470 2.570 ;
        RECT  3.010 3.440 3.250 3.840 ;
        RECT  3.210 1.550 3.230 1.790 ;
        RECT  2.970 1.390 3.210 1.790 ;
        RECT  2.950 2.870 3.190 3.110 ;
        RECT  2.430 3.440 3.010 3.680 ;
        RECT  2.710 2.070 2.950 3.110 ;
        RECT  2.690 2.070 2.710 2.310 ;
        RECT  2.450 0.870 2.690 2.310 ;
        RECT  2.190 2.910 2.430 3.680 ;
        RECT  2.170 2.910 2.190 3.310 ;
        RECT  1.930 1.390 2.170 3.310 ;
        RECT  1.840 2.910 1.930 3.310 ;
        RECT  1.670 3.650 1.910 4.360 ;
        RECT  1.470 3.650 1.670 3.890 ;
        RECT  1.470 2.010 1.650 2.410 ;
        RECT  1.230 1.180 1.470 3.890 ;
        RECT  0.570 1.180 1.230 1.420 ;
        RECT  0.170 3.490 1.230 3.890 ;
        RECT  0.170 1.020 0.570 1.420 ;
    END
END ADDFX4

MACRO ADDFX2
    CLASS CORE ;
    FOREIGN ADDFX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ ADDFXL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.610 3.130 14.730 4.110 ;
        RECT  14.720 2.390 14.730 2.650 ;
        RECT  14.610 0.820 14.730 1.950 ;
        RECT  14.730 0.820 14.970 4.110 ;
        RECT  14.970 2.390 14.980 2.650 ;
        RECT  14.970 3.130 15.010 4.110 ;
        RECT  14.970 0.820 15.010 1.950 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  13.080 2.890 13.240 3.290 ;
        RECT  13.080 0.730 13.240 1.710 ;
        RECT  13.240 0.730 13.480 3.290 ;
        RECT  13.480 2.390 13.660 2.650 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.970 1.960 10.010 2.200 ;
        RECT  10.100 2.950 10.130 3.210 ;
        RECT  10.010 1.960 10.130 2.400 ;
        RECT  10.130 1.960 10.370 3.360 ;
        RECT  10.370 2.950 10.620 3.360 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.220 2.090 ;
        RECT  0.220 1.830 0.460 2.420 ;
        RECT  0.460 2.010 0.700 2.420 ;
        RECT  0.700 2.010 0.810 2.410 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.280 2.320 5.260 2.720 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 4.480 1.390 5.440 ;
        RECT  1.390 4.640 9.920 5.440 ;
        RECT  9.920 3.840 9.930 5.440 ;
        RECT  9.930 3.640 10.330 5.440 ;
        RECT  10.330 3.840 10.340 5.440 ;
        RECT  10.340 4.640 13.850 5.440 ;
        RECT  13.850 4.090 14.250 5.440 ;
        RECT  14.250 4.640 15.180 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        RECT  0.990 -0.400 1.390 0.560 ;
        RECT  1.390 -0.400 4.880 0.400 ;
        RECT  4.880 -0.400 4.890 0.730 ;
        RECT  4.890 -0.400 5.290 0.850 ;
        RECT  5.290 -0.400 5.300 0.730 ;
        RECT  5.300 -0.400 10.570 0.400 ;
        RECT  10.570 -0.400 10.970 0.560 ;
        RECT  10.970 -0.400 13.840 0.400 ;
        RECT  13.840 -0.400 13.850 1.220 ;
        RECT  13.850 -0.400 14.250 1.710 ;
        RECT  14.250 -0.400 14.260 1.220 ;
        RECT  14.260 -0.400 15.180 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  14.260 2.180 14.360 2.580 ;
        RECT  14.020 2.180 14.260 3.810 ;
        RECT  13.520 3.570 14.020 3.810 ;
        RECT  13.280 3.570 13.520 4.130 ;
        RECT  11.980 3.890 13.280 4.130 ;
        RECT  12.560 0.710 12.800 3.590 ;
        RECT  12.340 0.710 12.560 1.100 ;
        RECT  12.340 3.190 12.560 3.590 ;
        RECT  10.330 0.860 12.340 1.100 ;
        RECT  11.850 3.200 11.980 4.130 ;
        RECT  11.850 1.430 11.930 1.830 ;
        RECT  11.740 1.430 11.850 4.130 ;
        RECT  11.610 1.430 11.740 3.600 ;
        RECT  11.530 1.430 11.610 1.830 ;
        RECT  11.580 3.200 11.610 3.600 ;
        RECT  11.520 1.510 11.530 1.750 ;
        RECT  10.900 1.430 11.140 3.600 ;
        RECT  10.650 1.430 10.900 1.830 ;
        RECT  9.850 1.430 10.650 1.670 ;
        RECT  10.090 0.680 10.330 1.100 ;
        RECT  6.610 0.680 10.090 0.920 ;
        RECT  9.610 1.200 9.850 1.670 ;
        RECT  9.460 2.320 9.650 2.720 ;
        RECT  7.210 1.200 9.610 1.440 ;
        RECT  9.450 2.310 9.460 3.280 ;
        RECT  9.370 2.310 9.450 3.480 ;
        RECT  9.130 1.720 9.370 3.480 ;
        RECT  9.050 2.310 9.130 3.480 ;
        RECT  9.040 2.310 9.050 3.280 ;
        RECT  8.370 1.720 8.610 4.360 ;
        RECT  8.090 3.960 8.370 4.360 ;
        RECT  7.850 1.950 8.090 3.410 ;
        RECT  7.730 1.950 7.850 2.190 ;
        RECT  7.450 3.170 7.850 3.410 ;
        RECT  7.490 1.720 7.730 2.190 ;
        RECT  7.500 2.480 7.570 2.880 ;
        RECT  7.210 2.470 7.500 2.880 ;
        RECT  7.290 3.170 7.450 3.570 ;
        RECT  7.050 3.170 7.290 4.360 ;
        RECT  6.970 1.200 7.210 2.880 ;
        RECT  5.820 4.050 7.050 4.360 ;
        RECT  6.690 2.640 6.970 2.880 ;
        RECT  5.870 1.930 6.690 2.330 ;
        RECT  6.530 2.640 6.690 3.510 ;
        RECT  6.370 0.680 6.610 1.590 ;
        RECT  6.450 2.640 6.530 3.770 ;
        RECT  6.290 3.110 6.450 3.770 ;
        RECT  6.210 1.130 6.370 1.590 ;
        RECT  3.770 3.530 6.290 3.770 ;
        RECT  4.610 1.130 6.210 1.370 ;
        RECT  5.870 3.010 5.930 3.250 ;
        RECT  5.630 1.650 5.870 3.250 ;
        RECT  1.910 4.120 5.820 4.360 ;
        RECT  4.090 1.650 5.630 1.890 ;
        RECT  4.050 3.010 5.630 3.250 ;
        RECT  4.370 0.870 4.610 1.370 ;
        RECT  2.690 0.870 4.370 1.110 ;
        RECT  3.850 1.390 4.090 1.890 ;
        RECT  3.530 2.330 3.770 3.770 ;
        RECT  3.470 2.330 3.530 2.570 ;
        RECT  3.230 1.550 3.470 2.570 ;
        RECT  3.010 3.440 3.250 3.840 ;
        RECT  3.210 1.550 3.230 1.790 ;
        RECT  2.970 1.390 3.210 1.790 ;
        RECT  2.950 2.870 3.190 3.110 ;
        RECT  2.430 3.440 3.010 3.680 ;
        RECT  2.710 2.070 2.950 3.110 ;
        RECT  2.690 2.070 2.710 2.310 ;
        RECT  2.450 0.870 2.690 2.310 ;
        RECT  2.190 2.910 2.430 3.680 ;
        RECT  2.170 2.910 2.190 3.310 ;
        RECT  1.930 1.390 2.170 3.310 ;
        RECT  1.840 2.910 1.930 3.310 ;
        RECT  1.670 3.650 1.910 4.360 ;
        RECT  1.470 3.650 1.670 3.890 ;
        RECT  1.470 2.010 1.650 2.410 ;
        RECT  1.230 1.180 1.470 3.890 ;
        RECT  0.570 1.180 1.230 1.420 ;
        RECT  0.170 3.490 1.230 3.890 ;
        RECT  0.170 1.020 0.570 1.420 ;
    END
END ADDFX2

MACRO ADDFX1
    CLASS CORE ;
    FOREIGN ADDFX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    LEQ ADDFXL ;
    SIZE 15.180 BY 5.040 ;
    SYMMETRY x y ;
    SITE umc6site ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  12.850 3.060 13.090 3.460 ;
        RECT  13.090 1.320 13.250 3.460 ;
        RECT  13.250 1.320 13.330 3.300 ;
        RECT  13.330 1.320 13.490 1.720 ;
        RECT  13.330 2.390 13.660 2.650 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER met1 ;
        RECT  14.370 2.970 14.730 3.370 ;
        RECT  14.720 2.390 14.730 2.650 ;
        RECT  14.610 1.340 14.730 1.980 ;
        RECT  14.730 1.340 14.770 3.370 ;
        RECT  14.770 1.340 14.970 3.290 ;
        RECT  14.970 2.390 14.980 2.650 ;
        RECT  14.970 1.340 15.010 1.980 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  9.970 1.960 10.010 2.200 ;
        RECT  10.010 1.960 10.150 2.400 ;
        RECT  10.150 1.960 10.390 4.350 ;
        RECT  10.390 3.950 10.630 4.350 ;
        RECT  10.630 4.060 11.020 4.340 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  0.200 1.830 0.210 2.090 ;
        RECT  0.210 1.830 0.460 2.420 ;
        RECT  0.460 2.010 0.570 2.420 ;
        RECT  0.570 2.010 0.810 2.410 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER met1 ;
        RECT  4.280 2.320 5.260 2.720 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 4.640 0.990 5.440 ;
        RECT  0.990 4.480 1.390 5.440 ;
        RECT  1.390 4.640 9.460 5.440 ;
        RECT  9.460 4.280 9.470 5.440 ;
        RECT  9.470 4.080 9.870 5.440 ;
        RECT  9.870 4.280 9.880 5.440 ;
        RECT  9.880 4.640 13.600 5.440 ;
        RECT  13.600 3.220 13.610 5.440 ;
        RECT  13.610 3.020 14.010 5.440 ;
        RECT  14.010 3.220 14.020 5.440 ;
        RECT  14.020 4.640 15.180 5.440 ;
        END
    END VDD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER met1 ;
        RECT  0.000 -0.400 0.990 0.400 ;
        RECT  0.990 -0.400 1.390 0.560 ;
        RECT  1.390 -0.400 4.880 0.400 ;
        RECT  4.880 -0.400 4.890 0.730 ;
        RECT  4.890 -0.400 5.290 0.850 ;
        RECT  5.290 -0.400 5.300 0.730 ;
        RECT  5.300 -0.400 10.570 0.400 ;
        RECT  10.570 -0.400 10.970 0.560 ;
        RECT  10.970 -0.400 13.840 0.400 ;
        RECT  13.840 -0.400 13.850 1.470 ;
        RECT  13.850 -0.400 14.250 1.670 ;
        RECT  14.250 -0.400 14.260 1.470 ;
        RECT  14.260 -0.400 15.180 0.400 ;
        END
    END GND
    OBS
        LAYER met1 ;
        RECT  12.930 3.850 13.330 4.250 ;
        RECT  11.750 3.870 12.930 4.110 ;
        RECT  12.510 0.710 12.760 1.110 ;
        RECT  12.270 0.710 12.510 3.590 ;
        RECT  10.330 0.870 12.270 1.110 ;
        RECT  12.110 3.190 12.270 3.590 ;
        RECT  11.750 1.430 11.910 1.830 ;
        RECT  11.510 1.430 11.750 4.110 ;
        RECT  11.350 3.200 11.510 3.600 ;
        RECT  10.710 1.430 10.950 3.510 ;
        RECT  9.850 1.430 10.710 1.670 ;
        RECT  10.670 3.110 10.710 3.510 ;
        RECT  10.090 0.680 10.330 1.110 ;
        RECT  6.610 0.680 10.090 0.920 ;
        RECT  9.610 1.200 9.850 1.670 ;
        RECT  9.650 2.520 9.660 3.410 ;
        RECT  9.370 2.320 9.650 3.610 ;
        RECT  7.200 1.200 9.610 1.440 ;
        RECT  9.250 1.720 9.370 3.610 ;
        RECT  9.240 1.720 9.250 3.410 ;
        RECT  9.130 1.720 9.240 2.640 ;
        RECT  8.370 1.720 8.610 4.360 ;
        RECT  8.090 3.960 8.370 4.360 ;
        RECT  7.850 1.880 8.090 3.430 ;
        RECT  7.730 1.880 7.850 2.120 ;
        RECT  7.450 3.190 7.850 3.430 ;
        RECT  7.490 1.720 7.730 2.120 ;
        RECT  7.430 2.510 7.570 2.910 ;
        RECT  7.290 3.190 7.450 3.590 ;
        RECT  7.200 2.500 7.430 2.910 ;
        RECT  7.050 3.190 7.290 4.360 ;
        RECT  6.960 1.200 7.200 2.910 ;
        RECT  5.820 4.050 7.050 4.360 ;
        RECT  6.690 2.670 6.960 2.910 ;
        RECT  6.530 2.670 6.690 3.510 ;
        RECT  5.870 1.930 6.680 2.330 ;
        RECT  6.370 0.680 6.610 1.590 ;
        RECT  6.450 2.670 6.530 3.770 ;
        RECT  6.290 3.110 6.450 3.770 ;
        RECT  6.210 1.130 6.370 1.590 ;
        RECT  3.770 3.530 6.290 3.770 ;
        RECT  4.610 1.130 6.210 1.370 ;
        RECT  5.870 3.010 5.930 3.250 ;
        RECT  5.630 1.650 5.870 3.250 ;
        RECT  1.910 4.120 5.820 4.360 ;
        RECT  4.090 1.650 5.630 1.890 ;
        RECT  4.050 3.010 5.630 3.250 ;
        RECT  4.370 0.870 4.610 1.370 ;
        RECT  2.690 0.870 4.370 1.110 ;
        RECT  3.850 1.390 4.090 1.890 ;
        RECT  3.530 2.330 3.770 3.770 ;
        RECT  3.470 2.330 3.530 2.570 ;
        RECT  3.230 1.550 3.470 2.570 ;
        RECT  3.010 3.440 3.250 3.840 ;
        RECT  3.210 1.550 3.230 1.790 ;
        RECT  2.970 1.390 3.210 1.790 ;
        RECT  2.950 2.870 3.190 3.110 ;
        RECT  2.430 3.440 3.010 3.680 ;
        RECT  2.710 2.070 2.950 3.110 ;
        RECT  2.690 2.070 2.710 2.310 ;
        RECT  2.450 0.870 2.690 2.310 ;
        RECT  2.190 2.910 2.430 3.680 ;
        RECT  2.170 2.910 2.190 3.310 ;
        RECT  1.930 1.390 2.170 3.310 ;
        RECT  1.840 2.910 1.930 3.310 ;
        RECT  1.670 3.650 1.910 4.360 ;
        RECT  1.470 3.650 1.670 3.890 ;
        RECT  1.470 2.010 1.650 2.410 ;
        RECT  1.230 1.180 1.470 3.890 ;
        RECT  0.570 1.180 1.230 1.420 ;
        RECT  0.170 3.490 1.230 3.890 ;
        RECT  0.170 1.020 0.570 1.420 ;
    END
END ADDFX1

END LIBRARY
