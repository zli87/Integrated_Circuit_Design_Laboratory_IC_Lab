module INST_MEM_2 #(parameter ID_WIDTH=4, ADDR_WIDTH=32, DATA_WIDTH=16) (
// Glbal Signal
  	  input clk,
  	  input rst_n,
// slave interface
      // axi write address channel
      // src master
      input wire [ID_WIDTH-1:0]     awid_s_inf,
      input wire [ADDR_WIDTH-1:0] awaddr_s_inf,
      input wire [2:0]            awsize_s_inf,
      input wire [1:0]           awburst_s_inf,
      input wire [7:0]             awlen_s_inf,
      input wire                 awvalid_s_inf,
      // src slave
      output reg                 awready_s_inf,
      // -----------------------------

      // axi write data channel
      // src master
      input wire [DATA_WIDTH-1:0]  wdata_s_inf,
      input wire                   wlast_s_inf,
      input wire                  wvalid_s_inf,
      // src slave
      output reg                  wready_s_inf,

      // axi write response channel
      // src slave
      output reg  [ID_WIDTH-1:0]     bid_s_inf,
      output reg  [1:0]            bresp_s_inf,
      output reg                  bvalid_s_inf,
      // src master
      input wire                  bready_s_inf,
      // -----------------------------

      // axi read address channel
      // src master
      input wire [ID_WIDTH-1:0]     arid_s_inf,
      input wire [ADDR_WIDTH-1:0] araddr_s_inf,
      input wire [7:0]             arlen_s_inf,
      input wire [2:0]            arsize_s_inf,
      input wire [1:0]           arburst_s_inf,
      input wire                 arvalid_s_inf,
      // src slave
      output reg                 arready_s_inf,
      // -----------------------------

      // axi read data channel
      // slave
      output reg [ID_WIDTH-1:0]      rid_s_inf,
      output reg [DATA_WIDTH-1:0]  rdata_s_inf,
      output reg [1:0]             rresp_s_inf,
      output reg                   rlast_s_inf,
      output reg                  rvalid_s_inf,
      // master
      input wire                  rready_s_inf
      // -----------------------------
);
// Modify your "dat" in this directory path to initialized DRAM Value

parameter DRAM_p_r = "../00_TESTBED/DRAM/inst_2_file.dat";
// Modify DRAM_R_LAT           for Initial Read Data Latency,
//        DRAM_W_LAT           for Initial Write Data Latency
//        MAX_WAIT_READY_CYCLE for control the Upperlimit time to wait Response Ready Signal
//
//        reg [7:0] DRMA_r [0:8*1024-1] is the storage element in this simulation model

parameter DRAM_R_LAT = 90, DRAM_W_LAT =100, MAX_WAIT_READY_CYCLE=300;
reg	[7:0]	DRAM_r	[0:8*1024-1];

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Mzdao78RXjm8lwxgPldSlw/cOH6+KDurO5M+QZXVfDKkWFrD2iBdFltvGAqcUup/
ncVyL77JS1ZLuAmEnuuaQsrhLbcwmWGP6ugIqfKnNFVk6rNCKHv7gBS8RTV0bTrv
oVFJO9GIc8PIKOE3IStBQVtVAOdeZZTVi263bODKHxV2gJm5Rbn2gQ==
//pragma protect end_key_block
//pragma protect digest_block
R38BjrdqTg43+wJLgrtrwZ9czcI=
//pragma protect end_digest_block
//pragma protect data_block
uMETIPbBee5WkjRjnYeo1HHtuk6PsydeRzO5qDvoSpFF5s5kXVk/0zf+MkCb7k/F
Nl70XyHtsNW/J10HjCtjPGjaFm7kIOdNhZ42n0BrxBH+Lbth3YT9gdb2COiAnAff
AEAriaoy2BOCTF/rJ2dV6e53pD4W+S22Ie93Nfg00QO0jGXHdnj43zrNNNS7lVZ9
lMOBnwKBaxMSwzARXbGE4Q427ATLWeFfWZXqNuMQLTxRpTxk+pXqjjE92p89RgjJ
80d3MFRmx2TVSFgTgt6Sn0Wz/41Nfjs/D6w3qILdK0xtb0CnKjRKKT6lmVyz3AOt
yTtZnqyAN8AvIgn8M+SJf7gDZyfRAWRGYVDRO8/tiIoZ/+w5/G0Q+0WmH+94SOus
JA9qXEqK5dXAkctfa5yrCHTokw2ios0A6JpqVqQ3Du4quUI9JdpFvx9H9B9LxN5T
iK9HdZJKWp4YNQgmIF62e3pFS2BuGQ+ciKqUwjRpBpO0zuePmzBiDOYtlufSh933
dolMuvlOn4wod9VfOiQQO3uAGcLFtUWoE2cCOSc4tEymimZQH71f1GlS4bIEOV31
zTUhgkQy+N3ZXJ6FWQvw2gm8kGk7l7HmytWLNcNMLvRy0PYkt50L6155fWDDsrhn
13M90C4HtnlohL5CrRvQ1TYxAKR37/3ZBYlECfXI2MAIfdmuTIFHHuq0cLSRHMlJ
k7urTKxA+cex6jSz2RvELw354tYD/Xo7vv2xCAQM4mnktvxYhyqeoEtYAB5vlaNM
u/47s06vw6XYxbTjV7KfvBPzDS/zTwOaH7dWTeC8uqJrb1A+T0eIsET5Vo7u0EGM
BBwQYpfn3nBeb3bbqZRIYTol5zVNBlIUDhJ3o8Rgfy0tZ33VzXOC9LtHVn8YQebi
Y3fBayxsA9Kjh6pgoZdpKhRsoHoLG+duq5PBDRi5N2Sfz8nufTghSZI5leb5Gf7J
Q5prhJyTfbBrymObxYKWD9aCJqr1wXdCJ6m6MFbrsYwjUO7es4jhhgFxOweX0wJ3
L8yUaK3Ns//C5J1KzS0Sz7OBYCzvHPTw7vmmpyFIjLntju2f+F4e8arSaiwR7L+/
dYkQ3TiT1FMOS1/FwqbQMuDSVJBvQ2Kw1APvaO3fAHQ2hvXL5y3BDq494Yw3JUzD
ldK6DF55Akjh5H6U1QGSoPCO3tlUTf+gNacb0bp7E/IFJBRdZLVhB4TZwEnqVC/T
4pizS702G6Yit8nhKKusDZGIWmxlQ/skRGHqrw0+G03zdDZ9dL9QllmnPIOSiECj
okbucC129ZYGt91gEg7pyWUKRL1kgVOJcYzHbbolx4/YCOIc0jvWcUtmAjSHO6yj
1/D/sSlCVzg8qo1K0AjbJY/vtTVeWvXMqtz48daaAanv6Sc3GcZWoJ9/wKr0Zhga
V1B9pFi4F8ghHne2Cf21LaC4wCYQzNTsteCVCw/lZoQ7rMX/JtKWGXFHeYIdeHdf
fCu0jF0MZdWgxO18517BAudobHRi3P5JkanVWeCCoMmuFsnpfp8vaWQ0o4my75sF
x3JWFec7rBwLJdXtuVhrNoAeO5DuGVGud98bHVRw12OQT+yatPUMh5XMi5Ifx/vz
k65qRjrinBckbCxFytgfZn/3VkDgCbs1VHImyjOlu6D/d6HVmDA4spmhPXTUyk0d
MSnZIe4nG3I5po/ut0S5MhNwKd8QA7/rc4kG4Gj/TJ/PNEjOWKFJ038Zcrr5eZ1m
Oiv/9h++vrf0dBiBK3eBsgrWwIylqHSP1KsvZpOUVJWsnsGUybOJ8bU4/9R95De6
R52p6gDPBuFVoZZNlU+Up8mlxq5JVr/MdvMZp5U7hObuGQcwfUHLg6M45ounN+im
lHMXR3thsggVTL0SnZtfB5DKQ61piZt7gf4SjQFanG0nHbFyDcljxRPMcbhIV5pV
Pu2Ps9/oGVM44RtIhSrP1Yt1yXAEq0PWAsOGc8o8kVe8cmCFDCD4zwuqDFKg72a5
Xbr8K3/a+JW5R2pidMj50bUP2ujaTxjM5KZ+mHz61LMivcGqdzActKJ3vwhPquCW
BiMJIR43ooneXlPomzsTUMlcRCuhZzQYVYB4G2UUhsszK4dcrqRvovHNLiLvOthE
7zJKpI8kdtsoWBpSSxhwt3I4yqxFEpsQ6yJFn6UMF2mtYpNLnUDyt/I8vUv145gi
3L8gInb0Z4EkP6x+v7KKlTyuP1S2UlBNZPYJHAh+v/LFoOBh8GK1F4E3XWIYJ7Nx
0B4r08BKsuupAHFHUMD9Xmm6wWHucmHEIkHnE3QQ7M2vnOt9tDz33QC6judmwWtf
1zorlAoFWunLvegeMgibzbXP3tjxyyBLmSBn6zhW+h0YIn7OmL/T23whY/lCLNUh
Cb9iamUK+NeFinAjj4OXAGMUd2a7ycz6i9meuzqqwYnklHBfQfIBIQEm98e/HCJo
54LbJzeEbjHj3oUTXxM68hNSWeo31iFAUM3nxn+yXav2V/CPYv2f1HPKdb1wveCH
F8bDBwzKh2rB3RAEA0+JV/lzhi6GVyxxGjWR1MN3ZCvBKK9AsONT6CmqkdiTykHY
Iz7Po0o+TpWjXEIH9pO/ZmdPJeyKuzF1O3/JHaxQRmCUjBIYoh+0pGmlkHovVCRX
kFcftlzDh8yww9Cab+JeB4t7BBLdJkeMdeA1vsJKwYxSrlgpzCwXQwZGwy8eFIR/
SEWbLCjDm3XCi4rA0qBEWv/waDkdJsomvw6OkI9u2hylhoqgUvp81H9W5gQM2WhR
lVCoB9mRK+FhX6m6148CleDOKlG4WQdoGN+Fpt4+3OrP6JYNBJbdP6nAkIfaMIW5
kSlonSeEfHCMr2ToyfQW+7fVM4HSernBfqKWLj+pGood0L47JKbdgiZUje6SZstd
+pof5mg0OusdrerbzoVcUgZsBJISpsIyYemfV1cOrx+aTD2uH2MRA65ziRxpjfjF
eR8qkhw3t09nFMZYkkghm65T7Zd7PgzA4ymPM4JH4ApM0a0U4/iUW7C+7Xh8pDAD
J+1p46gX0BHYMtx1UB6jMQVxAEfY8t60KhNFM2TuJBlTSqb+IDLruVPjHPKyadSi
PEtYijQNFHDnEKstFWTxleRVl7UYAPN1SKoJfzeRZRi//K9LrLpWaD2rWmSA/S1+
kKqSzFlbgbzvjrOtHeYtdzpjsZus2Oa87JjysJcGE8aH7kHjmVls7RfBljcez7oa
tucaSfX2rXNsYXzSjF1P+S+LOJKzEzGsNBfw6hcnRAJGpTdrW/tg/hzbDOARcSYL
hEkb7Jkf07hMRFn4WdPqNx62Imoa7bFWaaXDhTNb5AJXEiLgmcCalBaFoFhtSETy
jLl3K70kWMyi4WFV0ViQIYg0KZfYS0wia8fCQl94GYc8r93CpNFjLG82qUgtBuOE
PYFwOMazoVsmNMW/YcbJgILWi76H2LT+dyVHScMPGpX/1aFpzYGNl5jvQhwAzj1Y
9KlD9AQYPPNv0rbD0cbJINfssv1Sxm+J3cZ+KCYZPpb34ULVG49nEB2GZvJCF54Y
sUkJDIBQsLVAj7D1eVdtPlG8FfvFcow/2VsiweQiQOWGWMOnLePj1vM/rCblGXxn
ULQsH3XbIe6uVIsdzBdskIKGcM/zUXwT9Dl9CApdXC6TsHuqP8FzQWHDny01pPfm
uT3mvipM4uYxV/DJakLxNC50e1+x6aZYd6mPkH3Znto54aCca5Cm1AQixcWDeRdu
dVUuvoJ2/z7Em1VJfujYnV9Ve9oa+pZiqdWyBs4JmdFfWr3oCotQP0LVV2BuCAiF
EHo43CLHTw7FILGMQamdBpZSCnYV1djZvuzgxEIGV1qw3zRWbCoBlQwAv6qednIA
oycpbQfFK02KFulXbg8DjaXoJC1jZ8DdGX4vu9yFFALXHvdIrFOPYK6NJItexeeF
ZI7J6fBHQQwDf7PaAZ+W3FwpNJlfkDlFsNNuSiYZyv20SWN+VphHjDsqj5Mqtzps
UqJg69BC5euckvYXeWybu2Eod4k91WD27VQCtIhprulDFmhx9brP272dahEaNrQB
PHuvth1ByNOrf7ZKDvDqMiYQCHqaBAiEKE0IKhVD3AAxBo95XdG8yYfST/N0uT3x
PNdSosAmSNX/2y5+01t/7RLFbGF6c7XuK+eozXTJIrGtjSe3j/J5bHGJ6kGUwzq2
7trda2tayN9Ye0sO/dI9jApFejC1oY9nHWtIpeMRVhSsx6jQ8IteQoHuVS/l0VMB
2tLdCXxbSDCMHhXEEjKrLDMd08BGMQapjRks+JX84GTvk5o7pNyB7x8boj77ptN6
LitxjBGPDAotlfWoFH10ByT9Vx86zCAml8ltDq3NtdLnvaEfno3idMK9b/fV/zLK
S7joHK2E8uzrHfA5JwzfJdySU9KqY5pSt19algYhO3KwdcEzZRAYQsOrpiWF7hl6
zYSsNaYeLHquRg4Mdy1zbiUVC7p9vNaWt7azYO7+B2vveKhqLJKv+yX1EIrTTBpm
uL9Alq4alWRRIgkJgY284qxsbdKZmo3HJ6yNgG0KbrGxkje8Wcg/6fj2z1a50HDX
v5l+7gyZi1vhubZeB7ndUN5nZO7j8y52Fpyv0FAM3NMsZZz6bU3dgNUDnWyUNKPc
M8SIsqVAcVFQZ2qWvey3bTWgZcQu5GfHG91TiAwMdA4sWAZVPn+B/aYPZcZtXnbA
Kdi9l5YY8DLH8b7E6Wk1W//ptT/OiyDG9CtnvccAFiMVc1zdKplxxNbvV+XIsu3L
nLywl7WWNBu78ZVrYXl++bR4C4xwj2KUT8u/gWo6ZFQlw7/d/jmzz2Cw/5LbcjPq
Ka51mMOS2Gh1YCpLE37gMrELgOv8AMNpZ5qKOA5hnBDAq6Nd14+J+vXy2lfd2XVZ
APsMZtDa6vQwY6CqxwvZCHcL8YpJ3LG7nPE6wGF2qHQwtd6qNIja8yJdRlE9dMVx
fMPRIOMGlDJfC8SHb7vevlbt7Vz9kOI2kTgT7xTr5jvFWwpVV4rl1Z64+rD2+kg7
FPMEst549bIRqioyLDD4ksyms5BwfTpMdm+t9eY6qmdLgiRO36RAZvNDSFWo8XtJ
vyTezJ7mMH09Ncxm/0l/63WN5PY3zLtUhKpKxp/FY9m6hwTQ854AFhrKzAhiWqqo
1XMuw9R0g6GC83TG+lDTYYVo1VCLe6q/h0tS1J75Gw/sN7AC2dLzXTKq6kEGSvL3
pt5lnlHWadthN8KNBape4c4jqTzgn6hfVarPOLqWPox9YoyTa0Kl+HQhX31REcxg
ovs7+ynUxjTmj/5/hXc7R2NQg9MIe76zyjZ0QEHKbHX5pC4+QqxO3CxHZ+HyRccM
TrQnKzejZKavKOigcvQWOqjbn88BFRiOmQEH0ebQJk1Xe7llAoGkBY2Sa1rArQtL
F1LCPKuqw6+JrMi5lKf2qtbwQm7dVHMc+RpIKDAdU8KGhWRI5kGkGagBTAabSJkl
KgzWoIiX1GmA12/+/Lpc+5uthYIkUpAepsznRGDTP40CafYXdIKpCMRiAc1KqwC2
Xg2qWJh076uUkQFFH69XghjWnrbQaSbotv6T1x22o0JzVZeaFEc/ISv4khjs2A16
6tNizXmd28JUISKljYzSK6j4OLAvLv9qduI9IhF174JrBHrpqDu/f1ZMVJd/TNMx
+gePfC4BCGqhwYEQ3UgwQSQ7PKuIklI9G6/Hc0vmRqMUJoFxajKvi3squ8VO1+Nv
KGkqja9az0UpH2xDvdgWS7Ax35DZByt+EPDIB3o5pXJPx9d5kR4VE4iZ49QMKSTy
ueFeSyhH6DSmVHqHBp6FOvaxqlhEaTzGQIbguwwi6gOO5UC7LTCnX1eJ84u9EbjK
N2Ye3w19sTD+ZnMmdkrLPd+LjBQ5IXtwgWvFxK7MYRQrsuCo7j3KkHJL+PV2aOhe
/2wOOixrUOid2xVGeu9Ezaq+OiZsj+XYqwG2jq3CBk32wz3auyMNV3bSnG7ZbUJK
UZPDeDjLOqkUQCxF8cY3VyeTmqoODDKhRPG9FqDJWqM+1d6ICWaTfRBo9MeNJqCI
JyUEKHOO+eiy879jKXzqorl43bAa1kQx4z4sa3jdJT6DphEH5nPKbOtPitPCI7vs
HnfY8A1aOt8hW1/bgPsYQujHHBqZHhX3KfmoS6s44X/KXXFXMGqoeh/gOZnOGhq4
REbh6PPfI12qLRa4WH3i8HdVSaM/hmvLS7xAItiJyKJ3U+ZsvHsXJanYHfaT/N9k
C6hzVd7ozbWgqevKCNhUsfbiDa0BazYhhnqghugjgK6wAZiEFBpTH9PspXAO54vc
ieS5ckxGK1i39dPnUOMb23lsZTUpW6NQCPkI8VeCZZZE3AXfvGt/rAlCGyqmR/Hn
IIdF9JQeOHG0IeMXOIo8OjooXu9h8qQx4jDpTPhbA24maOA+vpDSu3tXTdX/x8WF
5qypKUGYEt3ErH7bpdulYTHrpuxIdLkthEn83uBvKgvNENazNFD+3ca3aTA638ks
9JjCdfTexF2phP/kDLqdKiVDzll1MPvKpj4Gk3MLQzbxEUipd2NyHtiG5Kh77PNH
rrWWMtEgFmZuzSRmmAvvNzC0CBgUo760LdEca7FqxJi0Sn7hmuOQd/1GJsmJJjDY
ccSHdhcwxo+s/LMQ3E5vEN9KCWEPX0RZCpkTDBUOG+TkaAusIR0y9QJ57aYfhmr3
2iOa7UKKQHQ2EwKaS1p0p0VsuJ+v98g/Ldn6pRw5IaN0u89lG12/rvgxTTVQN2Ib
enMWCB73XP0MIlQlJ2gaad0S9/KgvdCKfAIIRZ5lxoFsy91mxViPvI0LADFEguoC
LSnFnAaCz//az172YTWXpbtNIh2SNFpCDR7Pm/b2F67f7Nx/goLfiQG9WR4RkNC5
RwzR9JgRYZ+bMWtfO0l94JZEz2ZYT3S+nS3yWpP31y2v6S1qVtu50xxvLhJNuH8E
Ph2Zkc8CNaOc+q4ZS5L/zg8OSjUYh9tJKXK1ALYY0o3GtDkoUv0Usth95X/HMBA6
aH3sWVvpsa/gSgNlnjEs4BvdsNXX6sElF+QTLq9YV0OU7aOqZC7MHpQRyOBxp211
CDR+bEUB5pITaNo6SO0Q47LU4TZTsZKcW8y+BSNTVhBcfHW5beC6/LAlFODaASnr
DcVT1LvH683rBsE88GY79h9Hhg64zUtVbInaW4FSUl2bt0nnxUza741E2GrebnuM
PottHqTRB56uU9R0aYQUSq/A8Z8qaMJ5Bzdmz1eNPOIoJBfTUlgGC8ZYSkOrzN8v
WmC/HyICddUyLZNGLmL/F9754k3Hxy9O7ymjwYuFG8x4gN+6P7RiIEE4dwG7NOSU
AdUIMQVdakQEZvCuuTDF/d+MvwkcJ+mvQKiL1jcp3MzQLUWfnbQ1pzDytin9Yem8
ztLn0oDu1Z+AtQ4kX6jUFRPs+zpRPXQe6bhi7yN2pW2oIBCVtrjWR/exG57ERnnC
KPdRVLSLWCfLIA5w01koU8jLM4ywIubt0dL+FXEc+iPveQy7IfW+HEmfRdKsi7Rb
DqlyCaPjCMNYzMzVCBZsyh1ARDQjV2hAqX4gPF2UcOTnYhYyfdvt9tR3JCL1Goo8
eAVV+nhW4OaHgzN+po1C30XX8jcBgGzrH+RMZD6fLVXUR99ikEdKysvBUS6Nmmkv
3HQZcegkKUhL3ba4flLZpgdGk08g6SHljev90XlrDEAOYxAob0mOoHuKZiHC1CXd
PmXSVKSYFOJZx4vVtoxKkldcZgK2schvbDLyZg8pCF+ek12ZZER1L4IzTSNBhFyO
ClG5NOBHJ1yLfIWlL5Kxg/h3OwWO0YSggEugKJtn9+iiWOFS2Z6qLv830wLl0eDC
3XX2suZe9+pJvN62cLCeVv76lmLligURLvjMbkmze352u0+LpLnIMYPqZPC5Cf85
PYV98gOPp4Lfo+cJ96RCtBgK14lf0D7SJ6LKeJQ6J7pk+RSLme0+D8ppW7IEG32n
YUYdU8Qj/ovHLGAOV4dpR2laUDm/xcWBHyY+INHETv+W2JJbgbI0QxLr2uFn6nRd
jUib3rKfNpt0tJtSynvhJ4oDimJkDe2eRDyfuypdtYZwhRLXfan+RuDj+dJE5N/7
SgGh04RPJx5IPe3B0kpNV3WFj7jp6sOPOVPadf1mPzckhGTlP8+XcStc+Vb6aRXk
JkjTS6wc52luh3wAIGDtoOfZpTT6AMoO1J3CGKb0zXEweeMf0DAu9CML9+0Tve/A
USqodISoUA+2Q8TFCUR29ErVcmqCfRu6kQlGU5dsQ7mCb+HiiAyCkwMhhD4P+xzq
tMzUTppYSImtE+FaW+356n9bXO5KHi/aB5Pv1iDx8r8s9zYUwvmtdebPgBrP0Kzm
defb/cWG3x4IrelrwO2KGkXXDWWrZ0vhw9SypKIwXyfxSLdf6d3KySJLydqTxhhl
Lz/UnqZ3m7RFplpxPjXAdneLCpEgkZvhI5lWif2JOOFP2xRTuGBodSEMUVxm/2jO
SM4Y7u8S+VmEg1WmsbqzK4Jr9XJ4PjScl9IglK5PuDVypjjUs8FVf6/BgmCu7fKV
wIIiH3uqF/UNQK5yUfaG/sXmYIImQJeiHSGFzET9qBmLNzXGNET8d/j3q/3vPPiQ
UufrE854WaJCbBueQks2UDJV1wN/6m1DMV4OLU9Ol+v0KNNB2g0N8bkAH/VuJ3Zy
3ndv1N3t4WYI8CJO80V5idaiZqkBib62+GL+7swNdFTqxH+Hi9YKxQu6YdqLpif6
+kFVWwmdBRbNDJGDUVOdTTreoDRLxZ0iuwnm9m3Alw8DYlyWGj2ze8RaCfVP+nF8
R7NjzePfySIgtSZDEO6dDfoUzLIwJSJFGahi+zZJx17bgonmmMz4PzaGCYjV1h8S
y/0hx3NkG5VLgm0LB7irm3xNCrl3PnwlIgZG/DJNP2cGd8HzPwAniWyldvmuV4Y6
bWp/TqqQpa2yWgpTmNbuhvNn/AU4GkVpe2a0NcQ5Nd8QGZh6WCvY7WmfcoKLaKh0
IkB+RwJGS7jsqF9QaFnjsThqtSnw95/ptDr+IplX4Ib48MrYhZzdSfpGfsg9uMcV
bdMcDd5TpTsSUPIKdevq3jJwb1emqz6+FYr3yGxDaYFz8RyoLZFZIItu4axmGixT
ZhWuJz4zULZMwc4nCfxChlhuUPSBdFoOsRpFZu13gaaY+3HY0OjlKh8+drhC0Eto
5c0GpumBIqPIRXtobeus+XFE/lubCJkdwNwr1EbyRzbNrUyftnTgC1BDSzBE3+Rt
wXOcAraPXMonBkzaoDhS88iMgzNQPGZpFTPUneSFaXSSAHI9PRdnpv9YiR5G7trX
udszyetGdTtfMQW/+p74+1UGMx1tReTO8uPdjzffRz7k5J2wVfEQ9CVDzw1+mNY+
Si3YyDL4pJX3y3Wvw+LL6nG7EyKOUHxPajpGbBq5kRNr9VzYEIrdZMexTvtjb7vm
thpZN+n5i2eyI2lvRk2XAi1gHc1tbDAZdfRSoNP9r3uX0lZqJ98Z6XnbgJhpTjKx
SOyo4mH/MQgtTi9MVUi+DK9aMlAvX8F5E7iNpC5lmHVpFEXcmhnoy73KdckX2n0S
tsGlwUevPjE42Uly5jXI72ZWCjogapJqwygml/FVfq7x75j1MUPEUnr2hXlTTbAS
rY6pjXpfhDklrqKv5KtBHu5BjlBhYGs7t1ixLAJnVoDcH/czH1SObRCUwVp0oucV
x+ys2KJlMNWJG7lW77y/gIq420fr4WmGTzy3c360e/PiETjdLru0eGyws9TU/bW/
3ecJY035z+4qNjLa5xC1UchOBJWlAA9Cgd7T/JHH0fdnIXAomhfYrdH5zpuvIYVr
xOM9pgy285+vJcOVaazwLMeDsv35Jnp6slYkUr+Vl3LfrVV4tycDTAaWhiD25C7A
xcapulh+aaj70Fj0nCdHQ3efIFVAghsG9phIq9xWovHKOU5mjMF6zueZCpDTuJbl
4dhNh7vLVEWK3fXONsLNqUfb9KQ4ai0in/gc305mGnv/dNCSK72jpKBx7yszV3WM
iwJf5D9oZ8h9d4C35irlPk4LpwImQOchFVE3AI22RlYQR8KkKTHdYgKR59Obv9U+
7sb1NFfB5t2Kv3bI7kEMhrpT8b3S7bhrNTO9pH8KtsElWc0uthPWo6ZTkhxlFGoY
uGKqMsh5Qgg0aP9BzQtMQphX/qHlLmnQ6EE0CyBYGLz0ptQs5PAn7fPy7EIdIs7a
sZolbly+dEcGuz4QPKDQuDr2DnrkW8cBXDQANC4WWwjHrT5Y2cUsb7Z0G0nHwK51
BC8INO1KNj6mGezI0z6MN1/ZVP/bGAEJnSfcEUPbbJamxvGwz5q84ANbO1FtlgZL
Pdsb+Swd4I/p2VhQC/RN7ODlDKfqb+tZwjAiWudeQbYQ+Cemw7fMpn2V//KczmYG
HxLfshlOcsCffPAl9Jtg/nT79v7oKtpr7Z23bad11osuertDvrMoDi/glDLTfy3b
/46maifj+hjdI3MaO6AV/zoQdj3eX50aDgo58Sa1dkwkpbNYMclLWqGjgw/JfGjs
cHigfF8XUzRbKhbpXyfK6qD6+pXuH3u3LoFLPuk48fBnVWWuuooHfT4PVQc5cvLR
eKBPGV7Q+pWZfjfVQyovH9FamFRLQYa4Xucp1x6xIIx/L9mQjrCFcjRKQdT4gJWn
8LjFeqOqMP2qxFvURg2eQrMOg/X2csMz0a7mKyjS97i9NxDKfOEhBb41PqBTP/t/
t37eP+69nwhbCPPg3KWFEF6EnrFpdgetRAvSidXj726yEAdSETv7EF2Yk8XD77W0
UriFgvbh9AsV2IPiVqdNmLHA3xA3mhYJFus0BGFiVxMui1N4zRF96ti4RyehVS9E
AHBdecdWxeOG/fNbpEo2fNk9yrzRH/K+Sxze0Jy/B/EIHp43/qUTKuihgr6jClLJ
NB31c1A4h7lIXmgoBvADMk+2O+c/eA3frRYGBxEqn5FbU4ABrKhO62BrpAV1SVwX
KCTxIFl+KRbiHUth1AJ5zzLBPMcG1jEpiNgkB9Hf6XoIGK3iq2XrOchHB3VUxMA5
Xzhra2yEAaucGhZfiyRWPIKx/QaXUhBEdxJmPZZ+46nSkgyKUw3sWtXYacMmRvLm
bQK2qNpUNID1OVQqEWnvbBmxfnDI+ztc1W/mR7NdWlps4PRak4kx//9FPAScuaaG
h7mhvb0HKM+8I4s0rxOuxOJBOaqQf1stfprIesi0RRCjmVi8+vztUSt3wv5Uhk6Z
ZfVbPeW6QquFez1KT4b1tiB1qljfmiZtQ/rVQHLoSvEqQh+6LA5jXthaGPZYBG/R
zUsa2IU3NwK3Blv3/V5etxOM6KytwD9dZ9Fm0pVamMN9ZUMJYmPpbZ+yvk8tOCh+
JUo3U1NBf5mgwrbzFK39OL+IcAY5lsuxsBn0kjplHTUSXgrn9XWZ/ggD7Bb2iHQF
BKTR9xmC5zqbP4jpQpk4rSLqlDUbuN/ObZHsx4upACgZ/fALryv4iVG0XqQa4gvB
DE1QUPDmIaMFOkqwIt0cx2OZZpyfc+4Wmv2riynrE2cuSCyPurVUBvSsm2bjB61I
0vRA3zbbJByqhUv3SytMODwWJYmS5/U+no5qksX/QgY3oKgVoCnD4fk9fXwc6ysf
IeyGscZsl3rA4INxugJZDaqiWKwtfwQgjwNmB+ur6ovMjPzoelDrbN017I0XwIWi
x+x1L4xGRzzSLKNUptDOudEBFhwrqr85wt510JJlRTNKxggFYJ3Bp58eUk9OlCym
J0D3sSN4cSkVrmlwy9AWMLlsCXRdB+o8gbB/bqQwSEESOkMNzZNdPFVXdSY+0ZSI
QTqXzf1kcbFzcz9VEhiw3eSSCwjZ/mPPzsACYC6ZclkxztOxsxBFdATIgScuTk7P
t/F/SHXXaWilyx51xVwni+usjhYhWDCJX5Vd1loHeLWzTYWjHW7p/HgbPQpo9S9/
Kzy/AEsrGwZxawdj58KhUgPxy0UQ6KfVDbg4tG/c0ALTxeuQFnarOdbk+ZGbQCc6
CktyhEUAU20Gb0DBu1cV3LNy9BptxmlsFpRYk+coIg4aBa+VY171RicDL37WYghC
RushMtcJraXHdrIUFeaZnH6tbT2HMtZ4mGMFgbVt3IJ9vYfPyxKRAP1UfgMJ0Fan
bZeSpMGIdGjAWSOg725sHbvsE863R4yw+okmY/lv/YMFHi+DE0ZNMNvlq03rK5OI
KwrWreZWOEUNmIxYLq1wpHlTFbIcwQ+mCuq6zvNTgTr15pGq60fLSe9FEBU1ni6O
UUSjIn3T2uzB8y24QWSkriI/c76FhsZDYMMvi8C9LkbmlqrNHjtrPPXRgLyPHW+m
N1VGabXO6VTB13BMpe8ckg9XVAcffkBeHWRjRxb85T8RCHQHrXIpyDC8sZaDfaNu
hSEr5s2tFmL+tiyM3XqvrRBcYT78POknq/lvBT3f4nAr6sMFv0KAJFgLZmqmpmpH
rztF8P9BNImplN69MurDnSCVg4e5ORwgxsOyD/oSlN/wbkoZpnhZk3PLtFduCaRw
YSG5LJV6c3MF+2zbqzSmmnxnwhlt0ti42cfaduLijzNxSLu2DvgcNtf1ui4zlXLy
FBGFH3RK5brV8vz3HKFTzrfpDLGgkCk6MVTyNq2NrFnjrWXR+HwCfBt6YtfiLP8N
84mu8WgeE20a7ohvMHxisumi1E20Z4/8EG/uMbyqlPSKKDMttc2GjZdV7+/P7t8n
OCJDuCugtsJ4//JJ26QucD4ZZf+VStEwzcxE/KPDSUFIs1oDy6Vtvy/Bb+5vaViK
cYTNOo5cda4WUNyxLHValF19nKU2O+CDcHxLKEOhUUhVmg/9Xcz6LQZ7Kd64tWtW
vgW1earL/7/cw0cpdFO4DLogIIuY1Ha47JgIf8ZdQfO9wwIDyBybfgD3228wdQ5Y
hhMY6T23Qrt/XMYzfuAMunaJWhl3yyJkOiDfMEa1Bnja2MaIYb79ynRXvHMvt9aZ
ZwJRQ9KnRtnuyN8XBL+eTIOXjwbrqgxxYADn//GqoqAHBYohgGziiX9FKM2rYOWh
iYFd1gH0gSCQC61MRiU5F5s309KLymynwBNRGr1ToQnycfHKgsyRRpNDsJWO2May
PQZoP56rnJ8qhl4B9nwhaLBrk4RmrDIaPKzCjOy2odASmc2HESaDkp+I7hvSi6m4
3xgm4HpGHKs8y7UKIJc/eYmtL+DET5QyNF+1u2uzJBv5tXxqHpHJfzACoGUsXREV
iEhgi3smdhxCaNPz+lgf9LN1NYbeD+OSKolyxb6v49juikLYzUVsvGdPDVSKA/Gn
PKDMHG/n/PYJ98N3v+RnIroq/7PjqpK92rhbz0WN2IVjwW+gco/4wdzWsBL/mAx2
mocJhNezk2pw06/rFJgmGAbtDvNo7CwGaf/0525Ey04GGdSt1QE3KM0lqPMdDsQX
+D3NYoJduu/sra0pQIU55h94/RksE+lHmln8WRIBzWVL0QWVO90SwcBkThzPizBP
Ou3a8DUoX5LdN6Vo7z6dL3AKfjET9FEkmEus0pCgYYQTAcPR2A7zhVLeYLYps34V
VreHEpvQ3lpR64ZtL0PP9vePgxLg35Sv5Sy/nFc47VmvMxAa+Xix8/V9H3l1xe0d
GBaV1A1ioU2zslnTHe8/mfQinCVjJ6okynsZdlahAMQwG7sQvIR4sKfzpaFZW7r2
TAxJIh1ZO9JJAY7PD709kkh+v/Iw0dD6n/kOO17AA03q+HRJ0IVwc/oKUYBIkJbs
m0T8w0vadM0GuZPjhvZ1zUz8Kf481JVh9zKmldg94TkHPwnZJ0V8gVdJmz2YwnUR
pgRFvwCRf5SxRytijxc+6tyaTGn8z3d9+DHDPenQZONdxUUUCufx1QtefoieIWP5
t5thSQUzr/8VylRjlQ0QP0aJ6/6/t26BPxCYN8gmL1MA9oVps6ZX2xAms8r/XSwX
E4QChX+kyGIKbQgpxS09ttBKLBQx46B27aNgOFYjcPN/+0odW8RSzSKPYJ+I4LPg
5KT6TFfBxTJznUF6dP/JqvVKsL3aJXyj7XdMlggqrA0RMAaHg5bw7mqZ/IodMvXx
y6eE8EOH2zj8CnzsXH8/FcTFvAY+VYoYqX09G8HAiCWDgYizvxQBsN57yE3soGLa
dkbIsxSLJJY2b6bWFuL5bxj2oQZzdTsFp8rmXLUGfYrDaAn8jZPtRvaUee2VCG5i
RtvMpXNKE311uqx9u17PLTTY2bHE8vd00ewjDNvevj09XZYezuSmWtiolWwYBQF0
1xdbNWduIO6VzbvaFHfandltmlRaHwL9gjI7BBHkRgQhv+2Pd03Nssr3H8FtGLnQ
KQSWjbuz/bLjQIcLT/JWwKv5GhpzX2EQ8ryRaSijJKp/8xXIVQIF5x7MspT+KVdx
0dDJhANhlHt4nMHTtcp5T38XfIUBLbJTsMS3P8au5XpWONQn7arvE3mRnLt+YVNc
yYuA2aQQpEWEVUpf8EAjiT6ZqqDJ392qCdOv12TASdIfoyY505cKGph3U1JdbQTZ
5Vy+4E3h1Tt8nBS0kCtTEzbb7Vg+D9nqj2bojChsrY7st1exT+6L0KyU8zZkzkvd
sVsgQIw3DbrGgN29YBnb8M07vmj+Udf6/22bn3j3m5hSYQ7vf6nuR+Kl3oUcn4s8
lhFrz95hMUJmOvkAvdr5ofepNE06HtywZ6OX5AUHXynufv9bXrfriG5y3T3e15EJ
ZoYNav4nCfwMGkWHur3fRsIXI0+SyQ4qOp67ABtsJWGgIo2iBsXd6x7O0D8tVsZa
B2ZVpIG9edpYO+Ta8hytpWHf4nYkejS8UNCJeh/V60Dr+DF/zTfA1awbjxo1LZ89
B2UbZMhJDhwk0EV+M/OK1zXmcebNUdCY98GG2DRyT4WRoNQT7WjLXK6hvU6tbVgx
cf5QRPO2iO0x55HlgK34hCDgNjlmozfwsw/tWDGxaMd2fKJodxmz+wOaQz1+pxvs
0kYyDRZRwpOWDTa95qP5mLwNlsC8n8VbgLQFsEB/NzAi+IIHwr2eb2OxbS5+SRkW
P9o1xh+NRWog+d9ZIqjAKwkTLs38ZxWp52On6ln5wztD2++R69cXSJ+WvyRvh4x2
hpeea19OTXQpKo4sam6TL2wTiio5TLi5bjy0IIiabJVOJo9nUtgMPHCGpIb3rZVY
N5k3Z2xFITQpLlE1fWsBU9T2/bcE0YFcYkgUUqF0GEkLdx+EfJaUSqFmrFsCM1rZ
Fkiox1SlCbnJtP5NC2Y5Noclpb9jPHcTKyzPyh35j0Wdc9wFgEE6WVHrsOXeJ5IW
Gd34psQheAa9nn3l/jBua3EMrRJN0tgWmxkEaMzg3Uuw1DqbcWKpBBoun2OszXWn
Dwys0sbuyK2okLVROZ+JG65bgn3DunTTvjan6qJS95eBA7Z8EGKlMAwylIa5ea1K
0y68kbmb/3oVswtiskpu5JMZ4GlGkJqxGHMFhC29G7ac7+n7VJJjAFb5RkmG+BMF
uo73uRGsAdeG2LBnG3vFHsa+5EsN+t/rbO4tTPVe5hG6z7fiGsNOGQko7kovEkcD
R4g1qUAWB6ixZhQuM3NLzkqAh3ZA9SBmWyqQkhBzm7NWTh+uS8fjqBL9Ta61eCnF
0zj+PIdepRWqDNsisJ/zyd2a5mWhOCFUq0TwriUMDEXGDEEtkRaeWhSWL5tD3HJ8
TOMZ9CvDRuvC5outUPm2CLLW0ytMd6y1effFT16ycTvb5sGmcM+SF3s+Y2d9VEwf
BC0VJibMThHDDsZ4WSDDQu5BjQBk4eyRHM79VSSfLGvlKiYLAO04ONFDGx5Jigiy
Li3Y94pRUpCBlWPO1fyaZiUwN9WyqjDsrEdVD66emLDW6KkwlT1GXPMCTRcWC/Gw
3z/5r4sDECxTSfNXvnRpfP0NSf3NWpq/V7reFv8wJpPeHTUmuEp4yrj2hfNTmRR/
NZIQvYc10KxXDuk+NBvFvAW864LOjMnWUMk0h78XgFlwar3qYw/5r37/ItuIUbY5
/+VXb5/HY0VBkvvt2CQ5Pge38z5giNCobh7dTnPJ40qcPOA+XO7MQOqpz+LgUneF
m3N1FKUDKkhfPgpgQaf9jJ0ww9Y8FkpiWq5vxLeAL1H0qDyzW1/U3wld9dGE/rTC
KbE58ynfxCryNyK3XMNiTMdX1QrfA4/ZayqHlVJVayXS+ExUTCzpwQF6sJZLlQsh
iuJuwi/qnwoKAcpWickeis2jBapBab9DBwgjJyW/yJry8Frn9rQPGJ3SqXgr+F/u
kJEd57N4j9fuTtLRDg9ThOqSPlFSvs5mkyB0a6A6wBj4nKgofNnOKkJjFsikBubW
bWKv6IenUvQI6CYaz6d6uqhj2vdUeZnN6xdjzyaxSGR3mmwCImDIGx5JDM2FNpyH
Kbpm16vAgMYzISdx2CmviPRgkU7jQJTkqTrNZPxPnAM314I+Ln1ny6EJyGRF/r7m
9/q6e0mhmEf5b55fvluntJrbBWUm3kxYBtlp+GPCLm4P6HP71iBLv73LsshB16q4
yn4BNmLWtwuifr0n4NAOFYol8duXZP6Pr8Kn0+VqofanYo/8EUPfa52KoTB+V9Pl
ChMaTTt26z5eSdsNj7Wi0o1OPoI8Hfq3R1JHWLUE3YEeSAm6UhdEDfXNU2HzB3JD
YEFWYory7/txAwrO7PgKZZ+TTAO8JEkziuf78AKj/y4y5WB0S7JriK2aun7Dp3Ah
RFH5hkuJ4YHJibZvAPu0JI7mWhJ6iQ3nSbqWCaTaIuGvShKS/4T+NJ2/9C5Vfxx0
hgvy0DcdN3fFlMdi5iuONrGlaWF8Ul3V06WnSyelrdg8tYJ0KVGDCkBo4/viERyp
IxPrevL8L7xcTG+CvhiZCfSqKXJUfahaAX+Z//an38RIWGiFwCl+AFCFIxXR6gpN
k6zCaCFCLY/2Z5VsVq9MpXfPTE3+m9gPGMIgE0nNChuQepYE/fI9/NrRkIgmr9nx
480RjhtiK5uNVkfthr1wcqxycZ+Krh2LbCEkBdQZZ3GSCU87qwgKq+61X51ja8IE
zDenf8tc9Jno76Rwn05Gp8ftOmeeGcZ2keUFCDcMHeZT7IpiyjlgnKLpKLf24ejm
GOUtkqIvY1QkWqU/FrrC1AHv5s3IWP/XYCA94h0u1d53EZmkfM23vjuDZdMRFdyh
477bMwiBBjQVqvREt3kpKLjXzQZZx6nzdff9bRTO+UHY3/GdzhvJC+wULzvl2PTw
ZrvSP3Vs3K8DRbe7Y34APH6r9KEOvvGCO9+/6YGGs9OcNF2UL1ShYxUFhPL4GMw7
GZfXvED/tkh5aofjE623TyCY8Z+EBsGCsRfKnjd5ZNQMii7vXbXXY2yvqQQ0raz7
f88XxhyOhLSKwJW0wC/8mE8LOqgWSqweu7B3KGYwWX9sR0EplBrLEB8aThrChqAR
qtxpBlzvOaAfUzwq1zPkwi2nYyZNXMx/NvZOsU3QSPWB+l2mF3hHz+Og55GWlWB/
7YPYWVwvLPY3B4kNUK1z7yOSFtT8PLbcVA94lDyMJUScHj+eJ3SpUeIw9uTMPY/3
h8fXcxS1r7K2+rRixn8wE6I6xN958J7BfPLW3UHwMUN++roveEScswKbgDr3h3c1
Py4np24ewxSJWHrrxAG/wILRW9IKByDmd+i/LNR0qcc4dJykvbxb1hNqV2M6eMGs
Nb5PrJlL7I3YQTttpqFXGEQ8vS7/WGXCOsy/f5ceflx41ecnNhXRaQ5cvrkpaVEh
WA+rvA3M33/s/SruHIjFNQxrrgo6GHCPWVDuHOZnGSQ6yrj64zQigieo6f83CJPe
EuaaVJwh58Da/t7MI2gQYs/aMT0++oNNbL9/F51ceMtQBxX+AOQ15i0avXOQTM7+
CwA1GbOk+eXUim+OD2L0ykglaKe71cAmmgoXpVgIjModEiBktvgPGFemYonBKwem
iRxK8E+prWxPCTszcD5MOcc3UOcpNbBq4dA6hl7s2VgzOTiZMn842b0MDgBkyKGA
Ywx64WRA16uFvpbP1bl8Ro42HLS6yMzy2XgWs1u3+w9qjdSNRUpx9jeT25FyM4+b
E5z/KZCO2ajjaQ+h6NGQklnpG1wRv2yoUs9PONHUdveIuOS0RDZoDi0vLq5rCkM4
ZLhWVd5UKUJiK+YMgFOp1PDCWakiQa2ERuU9gwGS0po6XPamPrjqYUSbDpH/sOkx
Frjz/BLk9PK2WvmFapkDfrmSgihCu+GAJ+BpR9w2Q8dsTBfbfo/EbMkRmskNKQuR
6AXFWMhuQCeOqv6/rq90/xnEvnSmmxBCbVE5kTy/yNZJAzSJSN7mSt08fNGXZ3G/
8nk64sK78pVfyxrGGeCFYf5FZqHN4rLn+GvaFL7BILfAgRhRXaWOgJXsg7S7DYl/
ISUd6H9GDUG8TPaQXlreRFTDtO22cUAOEPZ3y4CgIREPQs6pujlP+R2ASIgsUyhX
/Mnnlm5i0akCPrHf6CfNx4Mr3vn2s9aXK+rCxt1L4rudHf0O/W1/1JrCjgdBe+tU
yBv0MoMSjyEJib5XuxeRwRD8stsSKto3Tag2063sh1tWN4hpwZmaxoDbRFIhGUdK
c5tAB6de9bV8tRfjUjY85oIQskTQ678DloRqNMtkKnOcYtzZqMfp35axcISUPTlo
+h+Ur6pqZXG8Xku6uc9T2v7Si8GA0Iaxd54MMnBHDP6maMNR84Mv6pxf2hHhJSt0
HW4jG7Yynhey8S6DaifrPUlyoyiYQ16pbKSCXmfjYZd+MpTv9FkBe+hvaJOerDAS
AVs7vPehsl3ssVMUS414I6Tedmoa38qFUPanaqhMtqoXaaVfXIFpJMQMJ/YLnqJ+
Sh2pVC/R9JyywYI4cy0uKthA97IcXC3nFt5A7ztFLqJYEFG09AtKI8R3BDAfnblp
D7tHMxTD1/UlNCk3PGoRfcEXaT1IGItIMmZv8C4y8XkRAxB3Su1WUmafme5Etfq3
AffU7o72QzZ7cjAcF3xvNHeUMpe17tipMxVosf/99CoRiAnQYqqEfmR8RmXhutmY
pFzFBnrNgkgLcfqYH8uve8UYnESVm7ZoWRSa/yCqzX3n7K9fhhVb7b/m3sD/eSRz
sCvnXZfmEjB6i+keveEiOvTY+UyMFdA4txFRqRn1QLjeUsETScqv0TjkIx7Yqqct
2NcLpE4MhjaVUCtiIL1V/pKSA1KQBB4+uP99AqQSgNeFHPKVL14ak/BB4zefvwG6
GCSkwWvy1VP2ZNemP1amJN3eqIYg4yrf7hnC9OqLzd28vv04oIK/QWdtmVYLTqoO
pq2D0ggyzCiep/rExtaQF9JPjTpYtycQ1O40H4nWU2o+NCivFlsOBOTGzVbW77UG
rsocMRdEcmebVT7CNFYennL4K5+aGPTJGHFzZYJwM3dv86dEJV5YzJ42h/shutiQ
bJUkJO0e+XGG8T5qLbfvKrLfow/5pjY1VXkrg+I+pRzev0Er/7VQKf4Jqph+xpAg
l9xDFORjY5QxOaqsK2e1/9n5YWQaS7pK9/CdUPQeqzaX48/oG43ycYK1gpKHBkvz
xHB0AuGQC0lHhDQxTEhIFBUizSuJGJuk1KqBJY4N/fn58+mY/nipH7YqYuAP+wgk
p94keUTY9iW7v7+I2/HDuQKK5mKgVhBZXbcTLsBd25rhNscQWIAMYxj9XqLp5vJn
tSsuuTffgSIwyDkjBVA5lyK76o79Z/7+KVps9fwGUILcvtEgwpnfkLPBPfHih2Y5
DGtHDSd/JDPo4jGKZmgEu3Z0OYNMD6yudt8AZqROoXE8ykAX91mGyyMH3ekOxzkn
7QTAK3dex1LYEcHtyIMzoixf06G35A9BtRRSonABKTG3+9qoekn2pO7E5OuN1pMx
ExaASExj+C7EwK8kX96225IZUMXIMKIXbWzqq+kXM0M=
//pragma protect end_data_block
//pragma protect digest_block
Ik78NQ2gA4p4lRGW+v2R/UhbqRY=
//pragma protect end_digest_block
//pragma protect end_protected
